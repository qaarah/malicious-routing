// Reading file 'aes.asc'..

module chip (input clk, input rst, output \d_out[6] , output \d_out[7] , output \d_out[5] , output \d_out[4] , output \d_out[3] , output \d_out[0] , output \d_out[2] , output \d_out[1] , output d_vld, input \d_in[7] , input \d_in[5] , input \d_in[6] , input \d_in[3] , input \d_in[0] , input \d_in[4] , input \d_in[1] , input \d_in[2] );

wire n1;
// (0, 0, 'glb_netwk_0')
// (2, 6, 'lutff_global/s_r')
// (2, 8, 'lutff_global/s_r')
// (4, 9, 'lutff_global/s_r')
// (6, 0, 'logic_op_tnr_6')
// (6, 1, 'neigh_op_rgt_6')
// (6, 2, 'lutff_global/s_r')
// (6, 2, 'neigh_op_bnr_6')
// (7, 0, 'fabout')
// (7, 0, 'local_g1_6')
// (7, 0, 'logic_op_top_6')
// (7, 1, 'lutff_6/out')
// (7, 2, 'neigh_op_bot_6')
// (8, 0, 'logic_op_tnl_6')
// (8, 1, 'neigh_op_lft_6')
// (8, 2, 'neigh_op_bnl_6')
// (11, 8, 'lutff_global/s_r')
// (12, 9, 'lutff_global/s_r')

reg n2 = 0;
// (0, 0, 'glb_netwk_1')
// (4, 10, 'lutff_global/cen')
// (4, 12, 'lutff_global/cen')
// (4, 14, 'neigh_op_tnr_2')
// (4, 15, 'neigh_op_rgt_2')
// (4, 16, 'neigh_op_bnr_2')
// (5, 12, 'lutff_global/cen')
// (5, 14, 'glb2local_3')
// (5, 14, 'local_g0_7')
// (5, 14, 'lutff_7/in_0')
// (5, 14, 'neigh_op_top_2')
// (5, 15, 'glb2local_1')
// (5, 15, 'local_g0_5')
// (5, 15, 'lutff_2/out')
// (5, 15, 'lutff_7/in_2')
// (5, 15, 'sp4_r_v_b_37')
// (5, 16, 'neigh_op_bot_2')
// (5, 16, 'sp4_r_v_b_24')
// (6, 11, 'lutff_global/cen')
// (6, 14, 'neigh_op_tnl_2')
// (6, 14, 'sp4_v_t_37')
// (6, 15, 'neigh_op_lft_2')
// (6, 15, 'sp4_v_b_37')
// (6, 16, 'neigh_op_bnl_2')
// (6, 16, 'sp4_v_b_24')
// (6, 17, 'span4_horz_r_2')
// (6, 17, 'span4_vert_13')
// (7, 12, 'glb2local_0')
// (7, 12, 'glb2local_1')
// (7, 12, 'local_g0_4')
// (7, 12, 'local_g0_5')
// (7, 12, 'lutff_0/in_3')
// (7, 12, 'lutff_4/in_3')
// (7, 12, 'lutff_5/in_3')
// (7, 12, 'lutff_7/in_3')
// (7, 17, 'fabout')
// (7, 17, 'local_g1_6')
// (7, 17, 'span4_horz_r_6')
// (8, 12, 'glb2local_0')
// (8, 12, 'local_g0_4')
// (8, 12, 'lutff_3/in_1')
// (8, 12, 'lutff_7/in_1')
// (8, 13, 'glb2local_0')
// (8, 13, 'local_g0_4')
// (8, 13, 'lutff_3/in_3')
// (8, 17, 'span4_horz_r_10')
// (9, 13, 'glb2local_3')
// (9, 13, 'local_g0_7')
// (9, 13, 'lutff_0/in_3')
// (9, 17, 'span4_horz_r_14')
// (10, 17, 'span4_horz_l_14')

wire n3;
// (0, 0, 'glb_netwk_2')
// (9, 13, 'lutff_global/s_r')
// (10, 11, 'neigh_op_tnr_5')
// (10, 12, 'neigh_op_rgt_5')
// (10, 12, 'sp4_r_v_b_42')
// (10, 13, 'neigh_op_bnr_5')
// (10, 13, 'sp4_r_v_b_31')
// (10, 14, 'sp4_r_v_b_18')
// (10, 15, 'sp4_r_v_b_7')
// (11, 11, 'neigh_op_top_5')
// (11, 11, 'sp4_h_r_0')
// (11, 11, 'sp4_v_t_42')
// (11, 12, 'lutff_5/out')
// (11, 12, 'sp4_v_b_42')
// (11, 13, 'lutff_global/s_r')
// (11, 13, 'neigh_op_bot_5')
// (11, 13, 'sp4_v_b_31')
// (11, 14, 'sp4_v_b_18')
// (11, 15, 'sp4_v_b_7')
// (12, 11, 'neigh_op_tnl_5')
// (12, 11, 'sp4_h_r_13')
// (12, 12, 'neigh_op_lft_5')
// (12, 13, 'neigh_op_bnl_5')
// (13, 7, 'span4_vert_t_14')
// (13, 8, 'span4_vert_b_14')
// (13, 9, 'fabout')
// (13, 9, 'local_g1_2')
// (13, 9, 'span4_vert_b_10')
// (13, 10, 'span4_vert_b_6')
// (13, 11, 'span4_horz_13')
// (13, 11, 'span4_vert_b_2')

wire n4;
// (0, 0, 'glb_netwk_4')
// (1, 12, 'lutff_global/s_r')
// (4, 4, 'lutff_global/s_r')
// (4, 6, 'lutff_global/s_r')
// (4, 13, 'glb2local_0')
// (4, 13, 'local_g0_4')
// (4, 13, 'lutff_7/in_3')
// (5, 11, 'lutff_global/s_r')
// (5, 14, 'neigh_op_tnr_4')
// (5, 14, 'sp4_r_v_b_37')
// (5, 15, 'neigh_op_rgt_4')
// (5, 15, 'sp4_r_v_b_24')
// (5, 16, 'neigh_op_bnr_4')
// (5, 16, 'sp4_r_v_b_13')
// (6, 13, 'sp4_v_t_37')
// (6, 14, 'neigh_op_top_4')
// (6, 14, 'sp4_v_b_37')
// (6, 15, 'lutff_4/out')
// (6, 15, 'sp4_v_b_24')
// (6, 16, 'neigh_op_bot_4')
// (6, 16, 'sp4_v_b_13')
// (6, 17, 'fabout')
// (6, 17, 'local_g1_0')
// (6, 17, 'span4_vert_0')
// (7, 9, 'lutff_global/s_r')
// (7, 14, 'neigh_op_tnl_4')
// (7, 15, 'neigh_op_lft_4')
// (7, 16, 'neigh_op_bnl_4')
// (11, 4, 'lutff_global/s_r')

wire clk;
// (0, 0, 'glb_netwk_6')
// (0, 4, 'span4_vert_t_14')
// (0, 5, 'span4_vert_b_14')
// (0, 6, 'span4_vert_b_10')
// (0, 7, 'span4_vert_b_6')
// (0, 8, 'fabout')
// (0, 8, 'io_1/D_IN_0')
// (0, 8, 'io_1/PAD')
// (0, 8, 'local_g1_2')
// (0, 8, 'span4_vert_b_2')
// (1, 7, 'neigh_op_tnl_2')
// (1, 7, 'neigh_op_tnl_6')
// (1, 8, 'neigh_op_lft_2')
// (1, 8, 'neigh_op_lft_6')
// (1, 9, 'neigh_op_bnl_2')
// (1, 9, 'neigh_op_bnl_6')
// (1, 12, 'lutff_global/clk')
// (2, 3, 'lutff_global/clk')
// (2, 4, 'lutff_global/clk')
// (2, 5, 'lutff_global/clk')
// (2, 6, 'lutff_global/clk')
// (2, 7, 'lutff_global/clk')
// (2, 8, 'lutff_global/clk')
// (2, 10, 'lutff_global/clk')
// (2, 11, 'lutff_global/clk')
// (2, 12, 'lutff_global/clk')
// (2, 15, 'lutff_global/clk')
// (4, 3, 'lutff_global/clk')
// (4, 4, 'lutff_global/clk')
// (4, 6, 'lutff_global/clk')
// (4, 7, 'lutff_global/clk')
// (4, 8, 'lutff_global/clk')
// (4, 9, 'lutff_global/clk')
// (4, 10, 'lutff_global/clk')
// (4, 11, 'lutff_global/clk')
// (4, 12, 'lutff_global/clk')
// (4, 14, 'lutff_global/clk')
// (5, 3, 'lutff_global/clk')
// (5, 4, 'lutff_global/clk')
// (5, 5, 'lutff_global/clk')
// (5, 6, 'lutff_global/clk')
// (5, 7, 'lutff_global/clk')
// (5, 8, 'lutff_global/clk')
// (5, 9, 'lutff_global/clk')
// (5, 10, 'lutff_global/clk')
// (5, 11, 'lutff_global/clk')
// (5, 12, 'lutff_global/clk')
// (5, 15, 'lutff_global/clk')
// (6, 2, 'lutff_global/clk')
// (6, 3, 'lutff_global/clk')
// (6, 4, 'lutff_global/clk')
// (6, 5, 'lutff_global/clk')
// (6, 6, 'lutff_global/clk')
// (6, 7, 'lutff_global/clk')
// (6, 8, 'lutff_global/clk')
// (6, 9, 'lutff_global/clk')
// (6, 10, 'lutff_global/clk')
// (6, 11, 'lutff_global/clk')
// (7, 3, 'lutff_global/clk')
// (7, 4, 'lutff_global/clk')
// (7, 5, 'lutff_global/clk')
// (7, 6, 'lutff_global/clk')
// (7, 7, 'lutff_global/clk')
// (7, 8, 'lutff_global/clk')
// (7, 9, 'lutff_global/clk')
// (8, 3, 'lutff_global/clk')
// (8, 4, 'lutff_global/clk')
// (8, 5, 'lutff_global/clk')
// (8, 6, 'lutff_global/clk')
// (8, 7, 'lutff_global/clk')
// (8, 8, 'lutff_global/clk')
// (9, 3, 'lutff_global/clk')
// (9, 4, 'lutff_global/clk')
// (9, 5, 'lutff_global/clk')
// (9, 6, 'lutff_global/clk')
// (9, 7, 'lutff_global/clk')
// (9, 8, 'lutff_global/clk')
// (9, 9, 'lutff_global/clk')
// (9, 13, 'lutff_global/clk')
// (9, 14, 'lutff_global/clk')
// (11, 3, 'lutff_global/clk')
// (11, 4, 'lutff_global/clk')
// (11, 5, 'lutff_global/clk')
// (11, 6, 'lutff_global/clk')
// (11, 7, 'lutff_global/clk')
// (11, 8, 'lutff_global/clk')
// (11, 9, 'lutff_global/clk')
// (11, 10, 'lutff_global/clk')
// (11, 11, 'lutff_global/clk')
// (11, 13, 'lutff_global/clk')
// (12, 7, 'lutff_global/clk')
// (12, 9, 'lutff_global/clk')
// (12, 12, 'lutff_global/clk')

wire n6;
// (0, 3, 'span12_horz_13')
// (1, 3, 'sp12_h_r_14')
// (2, 3, 'sp12_h_r_17')
// (2, 6, 'sp4_h_r_11')
// (3, 3, 'sp12_h_r_18')
// (3, 6, 'sp4_h_r_22')
// (4, 3, 'local_g0_5')
// (4, 3, 'lutff_1/in_2')
// (4, 3, 'sp12_h_r_21')
// (4, 6, 'local_g2_3')
// (4, 6, 'lutff_7/in_0')
// (4, 6, 'sp4_h_r_35')
// (5, 3, 'sp12_h_r_22')
// (5, 3, 'sp4_r_v_b_46')
// (5, 4, 'local_g2_3')
// (5, 4, 'lutff_3/in_2')
// (5, 4, 'sp4_r_v_b_35')
// (5, 5, 'sp4_r_v_b_22')
// (5, 6, 'sp4_h_r_46')
// (5, 6, 'sp4_r_v_b_11')
// (5, 11, 'neigh_op_tnr_3')
// (5, 12, 'neigh_op_rgt_3')
// (5, 13, 'neigh_op_bnr_3')
// (6, 2, 'sp4_v_t_46')
// (6, 3, 'sp12_h_l_22')
// (6, 3, 'sp12_v_t_22')
// (6, 3, 'sp4_v_b_46')
// (6, 4, 'sp12_v_b_22')
// (6, 4, 'sp4_v_b_35')
// (6, 5, 'sp12_v_b_21')
// (6, 5, 'sp4_v_b_22')
// (6, 6, 'sp12_v_b_18')
// (6, 6, 'sp4_h_l_46')
// (6, 6, 'sp4_v_b_11')
// (6, 7, 'sp12_v_b_17')
// (6, 8, 'sp12_v_b_14')
// (6, 9, 'sp12_v_b_13')
// (6, 10, 'sp12_v_b_10')
// (6, 11, 'neigh_op_top_3')
// (6, 11, 'sp12_v_b_9')
// (6, 12, 'lutff_3/out')
// (6, 12, 'sp12_v_b_6')
// (6, 13, 'neigh_op_bot_3')
// (6, 13, 'sp12_v_b_5')
// (6, 14, 'sp12_v_b_2')
// (6, 15, 'sp12_v_b_1')
// (7, 11, 'neigh_op_tnl_3')
// (7, 12, 'neigh_op_lft_3')
// (7, 13, 'neigh_op_bnl_3')

reg n7 = 0;
// (0, 3, 'span12_horz_3')
// (1, 3, 'sp12_h_r_4')
// (2, 3, 'sp12_h_r_7')
// (3, 3, 'sp12_h_r_8')
// (4, 3, 'sp12_h_r_11')
// (4, 3, 'sp4_h_r_7')
// (5, 3, 'sp12_h_r_12')
// (5, 3, 'sp4_h_r_18')
// (5, 4, 'sp4_r_v_b_44')
// (5, 5, 'sp4_r_v_b_33')
// (5, 6, 'sp4_r_v_b_20')
// (5, 7, 'sp4_r_v_b_9')
// (6, 3, 'sp12_h_r_15')
// (6, 3, 'sp4_h_r_31')
// (6, 3, 'sp4_h_r_9')
// (6, 3, 'sp4_v_t_44')
// (6, 4, 'sp4_v_b_44')
// (6, 5, 'local_g2_1')
// (6, 5, 'lutff_3/in_2')
// (6, 5, 'sp4_v_b_33')
// (6, 6, 'sp4_v_b_20')
// (6, 7, 'local_g0_1')
// (6, 7, 'local_g1_1')
// (6, 7, 'lutff_0/in_2')
// (6, 7, 'lutff_1/in_2')
// (6, 7, 'lutff_2/in_2')
// (6, 7, 'lutff_3/in_3')
// (6, 7, 'sp4_h_r_9')
// (6, 7, 'sp4_v_b_9')
// (7, 1, 'sp4_r_v_b_25')
// (7, 2, 'sp4_r_v_b_12')
// (7, 3, 'local_g0_0')
// (7, 3, 'lutff_2/in_2')
// (7, 3, 'sp12_h_r_16')
// (7, 3, 'sp4_h_r_20')
// (7, 3, 'sp4_h_r_42')
// (7, 3, 'sp4_r_v_b_1')
// (7, 4, 'local_g2_4')
// (7, 4, 'local_g2_5')
// (7, 4, 'lutff_0/in_2')
// (7, 4, 'lutff_1/in_2')
// (7, 4, 'lutff_5/in_3')
// (7, 4, 'sp4_r_v_b_36')
// (7, 4, 'sp4_r_v_b_37')
// (7, 5, 'local_g0_0')
// (7, 5, 'local_g1_0')
// (7, 5, 'lutff_0/in_2')
// (7, 5, 'lutff_1/in_2')
// (7, 5, 'lutff_2/in_3')
// (7, 5, 'sp4_r_v_b_24')
// (7, 5, 'sp4_r_v_b_25')
// (7, 6, 'local_g2_4')
// (7, 6, 'lutff_4/in_2')
// (7, 6, 'sp4_r_v_b_12')
// (7, 6, 'sp4_r_v_b_13')
// (7, 7, 'local_g0_4')
// (7, 7, 'local_g1_4')
// (7, 7, 'lutff_0/in_2')
// (7, 7, 'lutff_1/in_2')
// (7, 7, 'lutff_7/in_3')
// (7, 7, 'sp4_h_r_20')
// (7, 7, 'sp4_r_v_b_0')
// (7, 7, 'sp4_r_v_b_1')
// (8, 0, 'span4_vert_25')
// (8, 1, 'sp4_v_b_25')
// (8, 2, 'sp4_v_b_12')
// (8, 3, 'local_g0_3')
// (8, 3, 'local_g1_3')
// (8, 3, 'lutff_0/in_2')
// (8, 3, 'lutff_1/in_2')
// (8, 3, 'lutff_6/in_3')
// (8, 3, 'sp12_h_r_19')
// (8, 3, 'sp4_h_l_42')
// (8, 3, 'sp4_h_r_33')
// (8, 3, 'sp4_v_b_1')
// (8, 3, 'sp4_v_t_36')
// (8, 3, 'sp4_v_t_37')
// (8, 4, 'sp4_v_b_36')
// (8, 4, 'sp4_v_b_37')
// (8, 5, 'local_g3_0')
// (8, 5, 'lutff_5/in_2')
// (8, 5, 'lutff_6/in_3')
// (8, 5, 'sp4_v_b_24')
// (8, 5, 'sp4_v_b_25')
// (8, 6, 'local_g0_5')
// (8, 6, 'local_g1_5')
// (8, 6, 'lutff_1/in_2')
// (8, 6, 'lutff_2/in_2')
// (8, 6, 'sp4_v_b_12')
// (8, 6, 'sp4_v_b_13')
// (8, 7, 'sp4_h_r_33')
// (8, 7, 'sp4_v_b_0')
// (8, 7, 'sp4_v_b_1')
// (9, 3, 'local_g0_4')
// (9, 3, 'lutff_4/in_2')
// (9, 3, 'sp12_h_r_20')
// (9, 3, 'sp4_h_r_44')
// (9, 4, 'sp4_r_v_b_38')
// (9, 5, 'sp4_r_v_b_27')
// (9, 6, 'local_g2_6')
// (9, 6, 'lutff_0/in_2')
// (9, 6, 'lutff_3/in_3')
// (9, 6, 'lutff_6/in_2')
// (9, 6, 'sp4_r_v_b_14')
// (9, 7, 'local_g2_4')
// (9, 7, 'local_g3_4')
// (9, 7, 'lutff_1/in_2')
// (9, 7, 'lutff_2/in_2')
// (9, 7, 'lutff_3/in_2')
// (9, 7, 'lutff_5/in_3')
// (9, 7, 'sp4_h_r_44')
// (9, 7, 'sp4_r_v_b_3')
// (10, 3, 'sp12_h_r_23')
// (10, 3, 'sp4_h_l_44')
// (10, 3, 'sp4_v_t_38')
// (10, 4, 'sp4_v_b_38')
// (10, 5, 'sp4_v_b_27')
// (10, 6, 'sp4_v_b_14')
// (10, 7, 'sp4_h_l_44')
// (10, 7, 'sp4_v_b_3')
// (10, 10, 'neigh_op_tnr_4')
// (10, 11, 'neigh_op_rgt_4')
// (10, 12, 'neigh_op_bnr_4')
// (11, 3, 'sp12_h_l_23')
// (11, 3, 'sp12_v_t_23')
// (11, 4, 'sp12_v_b_23')
// (11, 5, 'local_g2_4')
// (11, 5, 'lutff_0/in_2')
// (11, 5, 'sp12_v_b_20')
// (11, 6, 'local_g3_3')
// (11, 6, 'lutff_0/in_2')
// (11, 6, 'sp12_v_b_19')
// (11, 7, 'sp12_v_b_16')
// (11, 8, 'sp12_v_b_15')
// (11, 9, 'sp12_v_b_12')
// (11, 10, 'neigh_op_top_4')
// (11, 10, 'sp12_v_b_11')
// (11, 11, 'lutff_4/out')
// (11, 11, 'sp12_v_b_8')
// (11, 12, 'neigh_op_bot_4')
// (11, 12, 'sp12_v_b_7')
// (11, 13, 'sp12_v_b_4')
// (11, 14, 'sp12_v_b_3')
// (11, 15, 'sp12_v_b_0')
// (12, 10, 'neigh_op_tnl_4')
// (12, 11, 'neigh_op_lft_4')
// (12, 12, 'neigh_op_bnl_4')

wire n8;
// (0, 3, 'span12_horz_8')
// (1, 3, 'sp12_h_r_11')
// (2, 3, 'sp12_h_r_12')
// (3, 3, 'sp12_h_r_15')
// (4, 2, 'sp4_r_v_b_40')
// (4, 3, 'sp12_h_r_16')
// (4, 3, 'sp4_r_v_b_29')
// (4, 4, 'sp4_r_v_b_16')
// (4, 5, 'sp4_r_v_b_5')
// (4, 6, 'sp4_r_v_b_39')
// (4, 7, 'sp4_r_v_b_26')
// (4, 8, 'sp4_r_v_b_15')
// (4, 9, 'sp4_r_v_b_2')
// (5, 1, 'sp4_v_t_40')
// (5, 2, 'sp4_v_b_40')
// (5, 3, 'sp12_h_r_19')
// (5, 3, 'sp4_v_b_29')
// (5, 4, 'local_g0_0')
// (5, 4, 'lutff_4/in_2')
// (5, 4, 'sp4_v_b_16')
// (5, 5, 'sp4_v_b_5')
// (5, 5, 'sp4_v_t_39')
// (5, 6, 'sp4_v_b_39')
// (5, 7, 'sp4_v_b_26')
// (5, 8, 'sp4_v_b_15')
// (5, 9, 'sp4_h_r_9')
// (5, 9, 'sp4_v_b_2')
// (6, 3, 'local_g1_4')
// (6, 3, 'lutff_4/in_3')
// (6, 3, 'lutff_5/in_2')
// (6, 3, 'sp12_h_r_20')
// (6, 9, 'local_g0_4')
// (6, 9, 'local_g1_4')
// (6, 9, 'lutff_3/in_3')
// (6, 9, 'lutff_4/in_3')
// (6, 9, 'lutff_5/in_3')
// (6, 9, 'sp4_h_r_20')
// (7, 3, 'sp12_h_r_23')
// (7, 8, 'neigh_op_tnr_6')
// (7, 9, 'neigh_op_rgt_6')
// (7, 9, 'sp4_h_r_33')
// (7, 10, 'neigh_op_bnr_6')
// (8, 3, 'sp12_h_l_23')
// (8, 3, 'sp12_v_t_23')
// (8, 4, 'sp12_v_b_23')
// (8, 5, 'sp12_v_b_20')
// (8, 6, 'sp12_v_b_19')
// (8, 7, 'sp12_v_b_16')
// (8, 8, 'neigh_op_top_6')
// (8, 8, 'sp12_v_b_15')
// (8, 9, 'lutff_6/out')
// (8, 9, 'sp12_v_b_12')
// (8, 9, 'sp4_h_r_44')
// (8, 10, 'neigh_op_bot_6')
// (8, 10, 'sp12_v_b_11')
// (8, 11, 'sp12_v_b_8')
// (8, 12, 'sp12_v_b_7')
// (8, 13, 'sp12_v_b_4')
// (8, 14, 'sp12_v_b_3')
// (8, 15, 'sp12_v_b_0')
// (9, 8, 'neigh_op_tnl_6')
// (9, 9, 'neigh_op_lft_6')
// (9, 9, 'sp4_h_l_44')
// (9, 10, 'neigh_op_bnl_6')

reg n9 = 0;
// (0, 4, 'span12_horz_1')
// (1, 4, 'sp12_h_r_2')
// (2, 4, 'sp12_h_r_5')
// (3, 4, 'sp12_h_r_6')
// (4, 3, 'neigh_op_tnr_1')
// (4, 4, 'neigh_op_rgt_1')
// (4, 4, 'sp12_h_r_9')
// (4, 5, 'neigh_op_bnr_1')
// (5, 3, 'neigh_op_top_1')
// (5, 4, 'local_g1_2')
// (5, 4, 'lutff_1/out')
// (5, 4, 'lutff_5/in_0')
// (5, 4, 'sp12_h_r_10')
// (5, 5, 'neigh_op_bot_1')
// (6, 3, 'neigh_op_tnl_1')
// (6, 4, 'neigh_op_lft_1')
// (6, 4, 'sp12_h_r_13')
// (6, 5, 'neigh_op_bnl_1')
// (7, 4, 'sp12_h_r_14')
// (8, 4, 'sp12_h_r_17')
// (9, 4, 'sp12_h_r_18')
// (10, 4, 'sp12_h_r_21')
// (11, 4, 'sp12_h_r_22')
// (12, 4, 'sp12_h_l_22')

wire n10;
// (0, 4, 'span12_horz_11')
// (0, 4, 'span4_horz_7')
// (1, 4, 'sp12_h_r_12')
// (1, 4, 'sp4_h_r_18')
// (2, 4, 'sp12_h_r_15')
// (2, 4, 'sp4_h_r_31')
// (3, 1, 'sp4_r_v_b_42')
// (3, 2, 'sp4_r_v_b_31')
// (3, 3, 'sp4_r_v_b_18')
// (3, 4, 'sp12_h_r_16')
// (3, 4, 'sp4_h_r_42')
// (3, 4, 'sp4_r_v_b_7')
// (4, 0, 'span4_vert_42')
// (4, 1, 'sp4_v_b_42')
// (4, 2, 'sp4_v_b_31')
// (4, 3, 'local_g0_2')
// (4, 3, 'lutff_1/in_3')
// (4, 3, 'sp4_v_b_18')
// (4, 4, 'sp12_h_r_19')
// (4, 4, 'sp4_h_l_42')
// (4, 4, 'sp4_v_b_7')
// (5, 4, 'sp12_h_r_20')
// (6, 3, 'local_g3_7')
// (6, 3, 'lutff_3/in_3')
// (6, 3, 'lutff_5/in_3')
// (6, 3, 'lutff_7/in_3')
// (6, 3, 'sp4_r_v_b_47')
// (6, 4, 'sp12_h_r_23')
// (6, 4, 'sp4_r_v_b_34')
// (6, 5, 'sp4_r_v_b_23')
// (6, 6, 'sp4_r_v_b_10')
// (6, 9, 'neigh_op_tnr_6')
// (6, 10, 'neigh_op_rgt_6')
// (6, 11, 'neigh_op_bnr_6')
// (7, 2, 'sp4_v_t_47')
// (7, 3, 'sp4_v_b_47')
// (7, 4, 'sp12_h_l_23')
// (7, 4, 'sp12_v_t_23')
// (7, 4, 'sp4_v_b_34')
// (7, 5, 'sp12_v_b_23')
// (7, 5, 'sp4_v_b_23')
// (7, 6, 'sp12_v_b_20')
// (7, 6, 'sp4_v_b_10')
// (7, 7, 'sp12_v_b_19')
// (7, 8, 'local_g3_0')
// (7, 8, 'lutff_6/in_3')
// (7, 8, 'sp12_v_b_16')
// (7, 9, 'local_g0_6')
// (7, 9, 'local_g1_6')
// (7, 9, 'lutff_0/in_3')
// (7, 9, 'lutff_3/in_3')
// (7, 9, 'neigh_op_top_6')
// (7, 9, 'sp12_v_b_15')
// (7, 10, 'lutff_6/out')
// (7, 10, 'sp12_v_b_12')
// (7, 11, 'neigh_op_bot_6')
// (7, 11, 'sp12_v_b_11')
// (7, 12, 'sp12_v_b_8')
// (7, 13, 'sp12_v_b_7')
// (7, 14, 'sp12_v_b_4')
// (7, 15, 'sp12_v_b_3')
// (7, 16, 'sp12_v_b_0')
// (8, 9, 'neigh_op_tnl_6')
// (8, 10, 'neigh_op_lft_6')
// (8, 11, 'neigh_op_bnl_6')

reg n11 = 0;
// (0, 4, 'span12_horz_8')
// (1, 3, 'neigh_op_tnr_2')
// (1, 4, 'neigh_op_rgt_2')
// (1, 4, 'sp12_h_r_11')
// (1, 5, 'neigh_op_bnr_2')
// (2, 3, 'neigh_op_top_2')
// (2, 4, 'lutff_2/out')
// (2, 4, 'sp12_h_r_12')
// (2, 5, 'neigh_op_bot_2')
// (3, 3, 'neigh_op_tnl_2')
// (3, 4, 'neigh_op_lft_2')
// (3, 4, 'sp12_h_r_15')
// (3, 5, 'neigh_op_bnl_2')
// (4, 4, 'sp12_h_r_16')
// (5, 4, 'local_g1_3')
// (5, 4, 'lutff_3/in_3')
// (5, 4, 'sp12_h_r_19')
// (6, 4, 'sp12_h_r_20')
// (7, 4, 'sp12_h_r_23')
// (8, 4, 'sp12_h_l_23')

reg n12 = 0;
// (0, 4, 'span4_horz_2')
// (1, 4, 'sp4_h_r_15')
// (2, 4, 'local_g2_2')
// (2, 4, 'lutff_2/in_0')
// (2, 4, 'sp4_h_r_26')
// (3, 1, 'sp4_r_v_b_44')
// (3, 2, 'neigh_op_tnr_2')
// (3, 2, 'sp4_r_v_b_33')
// (3, 3, 'neigh_op_rgt_2')
// (3, 3, 'sp4_r_v_b_20')
// (3, 4, 'neigh_op_bnr_2')
// (3, 4, 'sp4_h_r_39')
// (3, 4, 'sp4_r_v_b_9')
// (4, 0, 'span4_vert_44')
// (4, 1, 'sp4_v_b_44')
// (4, 2, 'neigh_op_top_2')
// (4, 2, 'sp4_v_b_33')
// (4, 3, 'lutff_2/out')
// (4, 3, 'sp4_v_b_20')
// (4, 4, 'neigh_op_bot_2')
// (4, 4, 'sp4_h_l_39')
// (4, 4, 'sp4_v_b_9')
// (5, 2, 'neigh_op_tnl_2')
// (5, 3, 'neigh_op_lft_2')
// (5, 4, 'neigh_op_bnl_2')

reg n13 = 0;
// (0, 6, 'span12_horz_12')
// (1, 5, 'neigh_op_tnr_4')
// (1, 6, 'neigh_op_rgt_4')
// (1, 6, 'sp12_h_r_15')
// (1, 7, 'neigh_op_bnr_4')
// (2, 5, 'neigh_op_top_4')
// (2, 6, 'lutff_4/out')
// (2, 6, 'sp12_h_r_16')
// (2, 7, 'neigh_op_bot_4')
// (3, 5, 'neigh_op_tnl_4')
// (3, 6, 'neigh_op_lft_4')
// (3, 6, 'sp12_h_r_19')
// (3, 7, 'neigh_op_bnl_4')
// (4, 6, 'sp12_h_r_20')
// (5, 6, 'local_g1_7')
// (5, 6, 'lutff_3/in_1')
// (5, 6, 'sp12_h_r_23')
// (6, 6, 'sp12_h_l_23')

reg n14 = 0;
// (0, 6, 'span12_horz_7')
// (1, 6, 'sp12_h_r_8')
// (2, 6, 'local_g1_3')
// (2, 6, 'lutff_4/in_0')
// (2, 6, 'sp12_h_r_11')
// (3, 6, 'sp12_h_r_12')
// (4, 5, 'neigh_op_tnr_4')
// (4, 6, 'neigh_op_rgt_4')
// (4, 6, 'sp12_h_r_15')
// (4, 7, 'neigh_op_bnr_4')
// (5, 5, 'neigh_op_top_4')
// (5, 6, 'local_g0_4')
// (5, 6, 'lutff_4/out')
// (5, 6, 'lutff_5/in_1')
// (5, 6, 'sp12_h_r_16')
// (5, 7, 'neigh_op_bot_4')
// (6, 5, 'neigh_op_tnl_4')
// (6, 6, 'neigh_op_lft_4')
// (6, 6, 'sp12_h_r_19')
// (6, 7, 'neigh_op_bnl_4')
// (7, 6, 'sp12_h_r_20')
// (8, 6, 'sp12_h_r_23')
// (9, 6, 'sp12_h_l_23')

reg n15 = 0;
// (0, 6, 'span4_horz_9')
// (1, 6, 'sp4_h_r_20')
// (2, 6, 'sp4_h_r_33')
// (3, 6, 'sp4_h_r_44')
// (4, 6, 'sp4_h_l_44')
// (4, 6, 'sp4_h_r_0')
// (4, 6, 'sp4_h_r_6')
// (4, 7, 'sp4_r_v_b_36')
// (4, 7, 'sp4_r_v_b_38')
// (4, 8, 'sp4_h_r_1')
// (4, 8, 'sp4_h_r_4')
// (4, 8, 'sp4_h_r_7')
// (4, 8, 'sp4_r_v_b_25')
// (4, 8, 'sp4_r_v_b_27')
// (4, 9, 'sp4_r_v_b_12')
// (4, 9, 'sp4_r_v_b_14')
// (4, 10, 'sp4_r_v_b_1')
// (4, 10, 'sp4_r_v_b_3')
// (5, 6, 'local_g0_3')
// (5, 6, 'local_g1_5')
// (5, 6, 'lutff_1/in_2')
// (5, 6, 'lutff_4/in_2')
// (5, 6, 'lutff_5/in_0')
// (5, 6, 'lutff_6/in_2')
// (5, 6, 'sp4_h_r_13')
// (5, 6, 'sp4_h_r_19')
// (5, 6, 'sp4_v_t_36')
// (5, 6, 'sp4_v_t_38')
// (5, 7, 'local_g2_4')
// (5, 7, 'lutff_2/in_2')
// (5, 7, 'lutff_4/in_2')
// (5, 7, 'sp4_v_b_36')
// (5, 7, 'sp4_v_b_38')
// (5, 8, 'local_g0_1')
// (5, 8, 'local_g0_4')
// (5, 8, 'lutff_5/in_0')
// (5, 8, 'lutff_7/in_1')
// (5, 8, 'sp4_h_r_12')
// (5, 8, 'sp4_h_r_17')
// (5, 8, 'sp4_h_r_18')
// (5, 8, 'sp4_v_b_25')
// (5, 8, 'sp4_v_b_27')
// (5, 9, 'local_g0_4')
// (5, 9, 'local_g1_6')
// (5, 9, 'lutff_2/in_2')
// (5, 9, 'lutff_3/in_2')
// (5, 9, 'lutff_4/in_2')
// (5, 9, 'lutff_7/in_1')
// (5, 9, 'sp4_v_b_12')
// (5, 9, 'sp4_v_b_14')
// (5, 10, 'sp4_h_r_3')
// (5, 10, 'sp4_h_r_8')
// (5, 10, 'sp4_v_b_1')
// (5, 10, 'sp4_v_b_3')
// (6, 3, 'local_g2_7')
// (6, 3, 'local_g3_1')
// (6, 3, 'lutff_3/in_2')
// (6, 3, 'lutff_4/in_2')
// (6, 3, 'lutff_5/in_0')
// (6, 3, 'lutff_7/in_2')
// (6, 3, 'sp4_r_v_b_39')
// (6, 3, 'sp4_r_v_b_41')
// (6, 4, 'sp4_r_v_b_26')
// (6, 4, 'sp4_r_v_b_28')
// (6, 5, 'sp4_r_v_b_15')
// (6, 5, 'sp4_r_v_b_17')
// (6, 6, 'sp4_h_r_24')
// (6, 6, 'sp4_h_r_30')
// (6, 6, 'sp4_r_v_b_2')
// (6, 6, 'sp4_r_v_b_4')
// (6, 7, 'sp4_r_v_b_37')
// (6, 7, 'sp4_r_v_b_45')
// (6, 8, 'local_g3_4')
// (6, 8, 'local_g3_7')
// (6, 8, 'lutff_1/in_2')
// (6, 8, 'lutff_2/in_2')
// (6, 8, 'sp4_h_r_25')
// (6, 8, 'sp4_h_r_28')
// (6, 8, 'sp4_h_r_31')
// (6, 8, 'sp4_r_v_b_24')
// (6, 8, 'sp4_r_v_b_32')
// (6, 9, 'local_g2_5')
// (6, 9, 'local_g3_5')
// (6, 9, 'lutff_2/in_2')
// (6, 9, 'lutff_3/in_2')
// (6, 9, 'lutff_4/in_2')
// (6, 9, 'lutff_5/in_0')
// (6, 9, 'sp4_r_v_b_13')
// (6, 9, 'sp4_r_v_b_21')
// (6, 10, 'sp4_h_r_14')
// (6, 10, 'sp4_h_r_21')
// (6, 10, 'sp4_r_v_b_0')
// (6, 10, 'sp4_r_v_b_8')
// (7, 2, 'sp4_v_t_39')
// (7, 2, 'sp4_v_t_41')
// (7, 3, 'sp4_v_b_39')
// (7, 3, 'sp4_v_b_41')
// (7, 4, 'sp4_v_b_26')
// (7, 4, 'sp4_v_b_28')
// (7, 5, 'sp4_r_v_b_36')
// (7, 5, 'sp4_r_v_b_47')
// (7, 5, 'sp4_v_b_15')
// (7, 5, 'sp4_v_b_17')
// (7, 6, 'sp4_h_r_2')
// (7, 6, 'sp4_h_r_37')
// (7, 6, 'sp4_h_r_43')
// (7, 6, 'sp4_r_v_b_25')
// (7, 6, 'sp4_r_v_b_34')
// (7, 6, 'sp4_v_b_2')
// (7, 6, 'sp4_v_b_4')
// (7, 6, 'sp4_v_t_37')
// (7, 6, 'sp4_v_t_45')
// (7, 7, 'sp4_r_v_b_12')
// (7, 7, 'sp4_r_v_b_23')
// (7, 7, 'sp4_v_b_37')
// (7, 7, 'sp4_v_b_45')
// (7, 8, 'local_g3_1')
// (7, 8, 'lutff_6/in_2')
// (7, 8, 'sp4_h_r_36')
// (7, 8, 'sp4_h_r_41')
// (7, 8, 'sp4_h_r_42')
// (7, 8, 'sp4_r_v_b_1')
// (7, 8, 'sp4_r_v_b_10')
// (7, 8, 'sp4_v_b_24')
// (7, 8, 'sp4_v_b_32')
// (7, 9, 'local_g2_4')
// (7, 9, 'lutff_4/in_0')
// (7, 9, 'sp4_r_v_b_36')
// (7, 9, 'sp4_v_b_13')
// (7, 9, 'sp4_v_b_21')
// (7, 10, 'sp4_h_r_27')
// (7, 10, 'sp4_h_r_32')
// (7, 10, 'sp4_r_v_b_25')
// (7, 10, 'sp4_v_b_0')
// (7, 10, 'sp4_v_b_8')
// (7, 11, 'sp4_r_v_b_12')
// (7, 12, 'sp4_r_v_b_1')
// (8, 4, 'sp4_v_t_36')
// (8, 4, 'sp4_v_t_47')
// (8, 5, 'sp4_v_b_36')
// (8, 5, 'sp4_v_b_47')
// (8, 6, 'sp4_h_l_37')
// (8, 6, 'sp4_h_l_43')
// (8, 6, 'sp4_h_r_15')
// (8, 6, 'sp4_h_r_3')
// (8, 6, 'sp4_v_b_25')
// (8, 6, 'sp4_v_b_34')
// (8, 7, 'local_g0_4')
// (8, 7, 'local_g0_7')
// (8, 7, 'lutff_1/in_2')
// (8, 7, 'lutff_2/in_2')
// (8, 7, 'lutff_3/in_0')
// (8, 7, 'lutff_7/in_2')
// (8, 7, 'sp4_v_b_12')
// (8, 7, 'sp4_v_b_23')
// (8, 8, 'sp4_h_l_36')
// (8, 8, 'sp4_h_l_41')
// (8, 8, 'sp4_h_l_42')
// (8, 8, 'sp4_h_r_1')
// (8, 8, 'sp4_v_b_1')
// (8, 8, 'sp4_v_b_10')
// (8, 8, 'sp4_v_t_36')
// (8, 9, 'sp4_v_b_36')
// (8, 10, 'sp4_h_r_38')
// (8, 10, 'sp4_h_r_45')
// (8, 10, 'sp4_v_b_25')
// (8, 11, 'sp4_v_b_12')
// (8, 12, 'sp4_v_b_1')
// (9, 6, 'sp4_h_r_14')
// (9, 6, 'sp4_h_r_26')
// (9, 8, 'sp4_h_r_12')
// (9, 10, 'sp4_h_l_38')
// (9, 10, 'sp4_h_l_45')
// (9, 10, 'sp4_h_r_0')
// (10, 6, 'sp4_h_r_27')
// (10, 6, 'sp4_h_r_39')
// (10, 7, 'sp4_r_v_b_45')
// (10, 8, 'sp4_h_r_25')
// (10, 8, 'sp4_r_v_b_32')
// (10, 9, 'neigh_op_tnr_4')
// (10, 9, 'sp4_r_v_b_21')
// (10, 10, 'neigh_op_rgt_4')
// (10, 10, 'sp4_h_r_13')
// (10, 10, 'sp4_r_v_b_8')
// (10, 11, 'neigh_op_bnr_4')
// (11, 6, 'sp4_h_l_39')
// (11, 6, 'sp4_h_r_38')
// (11, 6, 'sp4_v_t_45')
// (11, 7, 'sp4_r_v_b_44')
// (11, 7, 'sp4_v_b_45')
// (11, 8, 'sp4_h_r_36')
// (11, 8, 'sp4_r_v_b_33')
// (11, 8, 'sp4_v_b_32')
// (11, 9, 'local_g1_4')
// (11, 9, 'local_g2_4')
// (11, 9, 'lutff_4/in_2')
// (11, 9, 'lutff_5/in_2')
// (11, 9, 'lutff_6/in_0')
// (11, 9, 'lutff_7/in_2')
// (11, 9, 'neigh_op_top_4')
// (11, 9, 'sp4_r_v_b_20')
// (11, 9, 'sp4_r_v_b_36')
// (11, 9, 'sp4_v_b_21')
// (11, 10, 'lutff_4/out')
// (11, 10, 'sp4_h_r_24')
// (11, 10, 'sp4_r_v_b_25')
// (11, 10, 'sp4_r_v_b_9')
// (11, 10, 'sp4_v_b_8')
// (11, 11, 'neigh_op_bot_4')
// (11, 11, 'sp4_r_v_b_12')
// (11, 12, 'sp4_r_v_b_1')
// (12, 6, 'sp4_h_l_38')
// (12, 6, 'sp4_v_t_44')
// (12, 7, 'sp4_v_b_44')
// (12, 8, 'sp4_h_l_36')
// (12, 8, 'sp4_v_b_33')
// (12, 8, 'sp4_v_t_36')
// (12, 9, 'neigh_op_tnl_4')
// (12, 9, 'sp4_v_b_20')
// (12, 9, 'sp4_v_b_36')
// (12, 10, 'neigh_op_lft_4')
// (12, 10, 'sp4_h_r_37')
// (12, 10, 'sp4_v_b_25')
// (12, 10, 'sp4_v_b_9')
// (12, 11, 'neigh_op_bnl_4')
// (12, 11, 'sp4_v_b_12')
// (12, 12, 'sp4_v_b_1')
// (13, 10, 'span4_horz_37')

reg n16 = 0;
// (0, 7, 'span12_horz_0')
// (1, 7, 'sp12_h_r_3')
// (2, 7, 'local_g1_4')
// (2, 7, 'lutff_3/in_0')
// (2, 7, 'sp12_h_r_4')
// (3, 7, 'sp12_h_r_7')
// (4, 7, 'sp12_h_r_8')
// (5, 6, 'neigh_op_tnr_2')
// (5, 7, 'neigh_op_rgt_2')
// (5, 7, 'sp12_h_r_11')
// (5, 8, 'neigh_op_bnr_2')
// (6, 6, 'neigh_op_top_2')
// (6, 7, 'lutff_2/out')
// (6, 7, 'sp12_h_r_12')
// (6, 8, 'neigh_op_bot_2')
// (7, 6, 'neigh_op_tnl_2')
// (7, 7, 'neigh_op_lft_2')
// (7, 7, 'sp12_h_r_15')
// (7, 8, 'neigh_op_bnl_2')
// (8, 7, 'sp12_h_r_16')
// (9, 7, 'sp12_h_r_19')
// (10, 7, 'sp12_h_r_20')
// (11, 7, 'sp12_h_r_23')
// (12, 7, 'sp12_h_l_23')

reg n17 = 0;
// (0, 7, 'span12_horz_1')
// (1, 7, 'sp12_h_r_2')
// (2, 7, 'local_g1_5')
// (2, 7, 'lutff_2/in_0')
// (2, 7, 'sp12_h_r_5')
// (3, 7, 'sp12_h_r_6')
// (4, 6, 'neigh_op_tnr_1')
// (4, 7, 'neigh_op_rgt_1')
// (4, 7, 'sp12_h_r_9')
// (4, 8, 'neigh_op_bnr_1')
// (5, 6, 'neigh_op_top_1')
// (5, 7, 'lutff_1/out')
// (5, 7, 'sp12_h_r_10')
// (5, 8, 'neigh_op_bot_1')
// (6, 6, 'neigh_op_tnl_1')
// (6, 7, 'neigh_op_lft_1')
// (6, 7, 'sp12_h_r_13')
// (6, 8, 'neigh_op_bnl_1')
// (7, 7, 'sp12_h_r_14')
// (8, 7, 'sp12_h_r_17')
// (9, 7, 'sp12_h_r_18')
// (10, 7, 'sp12_h_r_21')
// (11, 7, 'sp12_h_r_22')
// (12, 7, 'sp12_h_l_22')

reg n18 = 0;
// (0, 7, 'span12_horz_10')
// (1, 6, 'neigh_op_tnr_3')
// (1, 7, 'neigh_op_rgt_3')
// (1, 7, 'sp12_h_r_13')
// (1, 8, 'neigh_op_bnr_3')
// (2, 6, 'neigh_op_top_3')
// (2, 7, 'lutff_3/out')
// (2, 7, 'sp12_h_r_14')
// (2, 8, 'neigh_op_bot_3')
// (3, 6, 'neigh_op_tnl_3')
// (3, 7, 'neigh_op_lft_3')
// (3, 7, 'sp12_h_r_17')
// (3, 8, 'neigh_op_bnl_3')
// (4, 7, 'sp12_h_r_18')
// (5, 7, 'local_g1_5')
// (5, 7, 'lutff_6/in_0')
// (5, 7, 'sp12_h_r_21')
// (6, 7, 'sp12_h_r_22')
// (7, 7, 'sp12_h_l_22')

reg n19 = 0;
// (0, 7, 'span12_horz_8')
// (1, 6, 'neigh_op_tnr_2')
// (1, 7, 'neigh_op_rgt_2')
// (1, 7, 'sp12_h_r_11')
// (1, 8, 'neigh_op_bnr_2')
// (2, 6, 'neigh_op_top_2')
// (2, 7, 'lutff_2/out')
// (2, 7, 'sp12_h_r_12')
// (2, 8, 'neigh_op_bot_2')
// (3, 6, 'neigh_op_tnl_2')
// (3, 7, 'neigh_op_lft_2')
// (3, 7, 'sp12_h_r_15')
// (3, 8, 'neigh_op_bnl_2')
// (4, 7, 'sp12_h_r_16')
// (5, 7, 'local_g0_3')
// (5, 7, 'lutff_3/in_0')
// (5, 7, 'sp12_h_r_19')
// (6, 7, 'sp12_h_r_20')
// (7, 7, 'sp12_h_r_23')
// (8, 7, 'sp12_h_l_23')

reg n20 = 0;
// (0, 8, 'span12_horz_0')
// (1, 8, 'sp12_h_r_3')
// (2, 8, 'local_g1_4')
// (2, 8, 'lutff_5/in_0')
// (2, 8, 'sp12_h_r_4')
// (3, 8, 'sp12_h_r_7')
// (4, 8, 'sp12_h_r_8')
// (5, 7, 'neigh_op_tnr_2')
// (5, 8, 'neigh_op_rgt_2')
// (5, 8, 'sp12_h_r_11')
// (5, 9, 'neigh_op_bnr_2')
// (6, 7, 'neigh_op_top_2')
// (6, 8, 'lutff_2/out')
// (6, 8, 'sp12_h_r_12')
// (6, 9, 'neigh_op_bot_2')
// (7, 7, 'neigh_op_tnl_2')
// (7, 8, 'local_g1_2')
// (7, 8, 'lutff_6/in_1')
// (7, 8, 'neigh_op_lft_2')
// (7, 8, 'sp12_h_r_15')
// (7, 9, 'neigh_op_bnl_2')
// (8, 8, 'sp12_h_r_16')
// (9, 8, 'sp12_h_r_19')
// (10, 8, 'sp12_h_r_20')
// (11, 8, 'sp12_h_r_23')
// (12, 8, 'sp12_h_l_23')

reg n21 = 0;
// (0, 8, 'span12_horz_13')
// (1, 8, 'sp12_h_r_14')
// (2, 8, 'local_g1_1')
// (2, 8, 'lutff_6/in_0')
// (2, 8, 'sp12_h_r_17')
// (3, 8, 'sp12_h_r_18')
// (4, 7, 'neigh_op_tnr_7')
// (4, 8, 'neigh_op_rgt_7')
// (4, 8, 'sp12_h_r_21')
// (4, 9, 'neigh_op_bnr_7')
// (5, 7, 'neigh_op_top_7')
// (5, 8, 'local_g1_7')
// (5, 8, 'lutff_5/in_1')
// (5, 8, 'lutff_7/out')
// (5, 8, 'sp12_h_r_22')
// (5, 9, 'neigh_op_bot_7')
// (6, 7, 'neigh_op_tnl_7')
// (6, 8, 'neigh_op_lft_7')
// (6, 8, 'sp12_h_l_22')
// (6, 9, 'neigh_op_bnl_7')

reg n22 = 0;
// (0, 8, 'span12_horz_2')
// (1, 8, 'sp12_h_r_5')
// (2, 8, 'local_g0_6')
// (2, 8, 'lutff_5/in_1')
// (2, 8, 'sp12_h_r_6')
// (3, 8, 'sp12_h_r_9')
// (4, 8, 'sp12_h_r_10')
// (5, 7, 'neigh_op_tnr_3')
// (5, 8, 'neigh_op_rgt_3')
// (5, 8, 'sp12_h_r_13')
// (5, 9, 'neigh_op_bnr_3')
// (6, 7, 'neigh_op_top_3')
// (6, 8, 'lutff_3/out')
// (6, 8, 'sp12_h_r_14')
// (6, 9, 'neigh_op_bot_3')
// (7, 7, 'neigh_op_tnl_3')
// (7, 8, 'neigh_op_lft_3')
// (7, 8, 'sp12_h_r_17')
// (7, 9, 'neigh_op_bnl_3')
// (8, 8, 'sp12_h_r_18')
// (9, 8, 'sp12_h_r_21')
// (10, 8, 'sp12_h_r_22')
// (11, 8, 'sp12_h_l_22')

reg n23 = 0;
// (0, 8, 'span12_horz_5')
// (1, 8, 'sp12_h_r_6')
// (2, 8, 'sp12_h_r_9')
// (3, 8, 'sp12_h_r_10')
// (4, 8, 'sp12_h_r_13')
// (5, 8, 'sp12_h_r_14')
// (6, 8, 'sp12_h_r_17')
// (7, 8, 'sp12_h_r_18')
// (8, 7, 'neigh_op_tnr_7')
// (8, 8, 'local_g0_5')
// (8, 8, 'lutff_6/in_3')
// (8, 8, 'neigh_op_rgt_7')
// (8, 8, 'sp12_h_r_21')
// (8, 9, 'neigh_op_bnr_7')
// (9, 7, 'neigh_op_top_7')
// (9, 8, 'lutff_7/out')
// (9, 8, 'sp12_h_r_22')
// (9, 9, 'neigh_op_bot_7')
// (10, 7, 'neigh_op_tnl_7')
// (10, 8, 'neigh_op_lft_7')
// (10, 8, 'sp12_h_l_22')
// (10, 9, 'neigh_op_bnl_7')

reg n24 = 0;
// (0, 9, 'span12_horz_0')
// (1, 9, 'sp12_h_r_3')
// (2, 9, 'sp12_h_r_4')
// (3, 9, 'sp12_h_r_7')
// (4, 9, 'local_g1_0')
// (4, 9, 'lutff_5/in_0')
// (4, 9, 'sp12_h_r_8')
// (5, 8, 'neigh_op_tnr_2')
// (5, 9, 'neigh_op_rgt_2')
// (5, 9, 'sp12_h_r_11')
// (5, 10, 'neigh_op_bnr_2')
// (6, 8, 'neigh_op_top_2')
// (6, 9, 'local_g0_2')
// (6, 9, 'lutff_2/out')
// (6, 9, 'lutff_5/in_1')
// (6, 9, 'sp12_h_r_12')
// (6, 10, 'neigh_op_bot_2')
// (7, 8, 'neigh_op_tnl_2')
// (7, 9, 'neigh_op_lft_2')
// (7, 9, 'sp12_h_r_15')
// (7, 10, 'neigh_op_bnl_2')
// (8, 9, 'sp12_h_r_16')
// (9, 9, 'sp12_h_r_19')
// (10, 9, 'sp12_h_r_20')
// (11, 9, 'sp12_h_r_23')
// (12, 9, 'sp12_h_l_23')

reg n25 = 0;
// (0, 9, 'span12_horz_10')
// (1, 9, 'sp12_h_r_13')
// (2, 9, 'sp12_h_r_14')
// (3, 8, 'neigh_op_tnr_5')
// (3, 9, 'neigh_op_rgt_5')
// (3, 9, 'sp12_h_r_17')
// (3, 10, 'neigh_op_bnr_5')
// (4, 8, 'neigh_op_top_5')
// (4, 9, 'lutff_5/out')
// (4, 9, 'sp12_h_r_18')
// (4, 10, 'neigh_op_bot_5')
// (5, 8, 'neigh_op_tnl_5')
// (5, 9, 'neigh_op_lft_5')
// (5, 9, 'sp12_h_r_21')
// (5, 10, 'neigh_op_bnl_5')
// (6, 9, 'local_g1_6')
// (6, 9, 'lutff_0/in_1')
// (6, 9, 'sp12_h_r_22')
// (7, 9, 'sp12_h_l_22')

reg n26 = 0;
// (0, 10, 'span12_horz_0')
// (1, 9, 'neigh_op_tnr_6')
// (1, 10, 'neigh_op_rgt_6')
// (1, 10, 'sp12_h_r_3')
// (1, 11, 'neigh_op_bnr_6')
// (2, 9, 'neigh_op_top_6')
// (2, 10, 'lutff_6/out')
// (2, 10, 'sp12_h_r_4')
// (2, 11, 'neigh_op_bot_6')
// (3, 9, 'neigh_op_tnl_6')
// (3, 10, 'neigh_op_lft_6')
// (3, 10, 'sp12_h_r_7')
// (3, 11, 'neigh_op_bnl_6')
// (4, 10, 'sp12_h_r_8')
// (5, 10, 'sp12_h_r_11')
// (5, 10, 'sp4_h_r_7')
// (6, 10, 'local_g0_2')
// (6, 10, 'lutff_4/in_0')
// (6, 10, 'sp12_h_r_12')
// (6, 10, 'sp4_h_r_18')
// (7, 10, 'sp12_h_r_15')
// (7, 10, 'sp4_h_r_31')
// (8, 10, 'sp12_h_r_16')
// (8, 10, 'sp4_h_r_42')
// (9, 10, 'sp12_h_r_19')
// (9, 10, 'sp4_h_l_42')
// (10, 10, 'sp12_h_r_20')
// (11, 10, 'sp12_h_r_23')
// (12, 10, 'sp12_h_l_23')

reg n27 = 0;
// (0, 11, 'logic_op_tnr_0')
// (0, 12, 'logic_op_rgt_0')
// (0, 13, 'logic_op_bnr_0')
// (1, 11, 'neigh_op_top_0')
// (1, 12, 'lutff_0/out')
// (1, 13, 'neigh_op_bot_0')
// (2, 11, 'neigh_op_tnl_0')
// (2, 12, 'local_g0_0')
// (2, 12, 'lutff_4/in_0')
// (2, 12, 'neigh_op_lft_0')
// (2, 13, 'neigh_op_bnl_0')

reg n28 = 0;
// (0, 11, 'span12_horz_0')
// (1, 10, 'neigh_op_tnr_6')
// (1, 11, 'neigh_op_rgt_6')
// (1, 11, 'sp12_h_r_3')
// (1, 12, 'neigh_op_bnr_6')
// (2, 10, 'neigh_op_top_6')
// (2, 11, 'lutff_6/out')
// (2, 11, 'sp12_h_r_4')
// (2, 12, 'neigh_op_bot_6')
// (3, 10, 'neigh_op_tnl_6')
// (3, 11, 'neigh_op_lft_6')
// (3, 11, 'sp12_h_r_7')
// (3, 12, 'neigh_op_bnl_6')
// (4, 11, 'local_g0_0')
// (4, 11, 'local_g1_0')
// (4, 11, 'lutff_0/in_2')
// (4, 11, 'lutff_3/in_0')
// (4, 11, 'sp12_h_r_8')
// (5, 11, 'sp12_h_r_11')
// (6, 11, 'sp12_h_r_12')
// (7, 11, 'sp12_h_r_15')
// (8, 11, 'sp12_h_r_16')
// (9, 11, 'sp12_h_r_19')
// (10, 11, 'sp12_h_r_20')
// (11, 11, 'sp12_h_r_23')
// (12, 11, 'sp12_h_l_23')

reg n29 = 0;
// (0, 11, 'span12_horz_3')
// (1, 11, 'sp12_h_r_4')
// (2, 11, 'sp12_h_r_7')
// (3, 11, 'sp12_h_r_8')
// (4, 11, 'sp12_h_r_11')
// (5, 11, 'sp12_h_r_12')
// (6, 11, 'local_g1_7')
// (6, 11, 'lutff_1/in_3')
// (6, 11, 'sp12_h_r_15')
// (7, 11, 'sp12_h_r_16')
// (8, 11, 'sp12_h_r_19')
// (9, 11, 'sp12_h_r_20')
// (10, 3, 'sp4_r_v_b_36')
// (10, 4, 'neigh_op_tnr_6')
// (10, 4, 'sp4_r_v_b_25')
// (10, 5, 'neigh_op_rgt_6')
// (10, 5, 'sp4_r_v_b_12')
// (10, 6, 'neigh_op_bnr_6')
// (10, 6, 'sp4_r_v_b_1')
// (10, 11, 'sp12_h_r_23')
// (11, 0, 'span12_vert_20')
// (11, 1, 'sp12_v_b_20')
// (11, 2, 'sp12_v_b_19')
// (11, 2, 'sp4_v_t_36')
// (11, 3, 'sp12_v_b_16')
// (11, 3, 'sp4_v_b_36')
// (11, 4, 'neigh_op_top_6')
// (11, 4, 'sp12_v_b_15')
// (11, 4, 'sp4_v_b_25')
// (11, 5, 'lutff_6/out')
// (11, 5, 'sp12_v_b_12')
// (11, 5, 'sp4_v_b_12')
// (11, 6, 'local_g0_1')
// (11, 6, 'lutff_1/in_0')
// (11, 6, 'neigh_op_bot_6')
// (11, 6, 'sp12_v_b_11')
// (11, 6, 'sp4_v_b_1')
// (11, 7, 'sp12_v_b_8')
// (11, 8, 'sp12_v_b_7')
// (11, 9, 'sp12_v_b_4')
// (11, 10, 'sp12_v_b_3')
// (11, 11, 'sp12_h_l_23')
// (11, 11, 'sp12_v_b_0')
// (12, 4, 'neigh_op_tnl_6')
// (12, 5, 'neigh_op_lft_6')
// (12, 6, 'neigh_op_bnl_6')

wire n30;
// (0, 11, 'span12_horz_8')
// (1, 10, 'neigh_op_tnr_2')
// (1, 11, 'neigh_op_rgt_2')
// (1, 11, 'sp12_h_r_11')
// (1, 12, 'neigh_op_bnr_2')
// (2, 10, 'neigh_op_top_2')
// (2, 11, 'lutff_2/out')
// (2, 11, 'sp12_h_r_12')
// (2, 12, 'neigh_op_bot_2')
// (3, 10, 'neigh_op_tnl_2')
// (3, 11, 'neigh_op_lft_2')
// (3, 11, 'sp12_h_r_15')
// (3, 12, 'neigh_op_bnl_2')
// (4, 11, 'sp12_h_r_16')
// (5, 11, 'sp12_h_r_19')
// (6, 11, 'local_g0_4')
// (6, 11, 'local_g1_4')
// (6, 11, 'lutff_2/in_2')
// (6, 11, 'lutff_4/in_3')
// (6, 11, 'sp12_h_r_20')
// (7, 11, 'sp12_h_r_23')
// (8, 11, 'sp12_h_l_23')

wire n31;
// (0, 12, 'span12_horz_6')
// (1, 11, 'neigh_op_tnr_1')
// (1, 12, 'neigh_op_rgt_1')
// (1, 12, 'sp12_h_r_9')
// (1, 13, 'neigh_op_bnr_1')
// (2, 11, 'neigh_op_top_1')
// (2, 12, 'lutff_1/out')
// (2, 12, 'sp12_h_r_10')
// (2, 13, 'neigh_op_bot_1')
// (3, 11, 'neigh_op_tnl_1')
// (3, 12, 'neigh_op_lft_1')
// (3, 12, 'sp12_h_r_13')
// (3, 13, 'neigh_op_bnl_1')
// (4, 12, 'local_g0_6')
// (4, 12, 'lutff_5/in_1')
// (4, 12, 'sp12_h_r_14')
// (5, 12, 'sp12_h_r_17')
// (6, 12, 'sp12_h_r_18')
// (7, 12, 'sp12_h_r_21')
// (8, 12, 'sp12_h_r_22')
// (9, 12, 'sp12_h_l_22')

reg n32 = 0;
// (0, 12, 'span12_horz_8')
// (1, 11, 'neigh_op_tnr_2')
// (1, 12, 'neigh_op_rgt_2')
// (1, 12, 'sp12_h_r_11')
// (1, 13, 'neigh_op_bnr_2')
// (2, 2, 'sp12_v_t_23')
// (2, 3, 'sp12_v_b_23')
// (2, 4, 'sp12_v_b_20')
// (2, 5, 'sp12_v_b_19')
// (2, 6, 'sp12_v_b_16')
// (2, 7, 'sp12_v_b_15')
// (2, 8, 'local_g2_4')
// (2, 8, 'lutff_5/in_3')
// (2, 8, 'sp12_v_b_12')
// (2, 9, 'sp12_v_b_11')
// (2, 9, 'sp4_r_v_b_40')
// (2, 10, 'sp12_v_b_8')
// (2, 10, 'sp4_r_v_b_29')
// (2, 11, 'neigh_op_top_2')
// (2, 11, 'sp12_v_b_7')
// (2, 11, 'sp4_r_v_b_16')
// (2, 12, 'lutff_2/out')
// (2, 12, 'sp12_h_r_12')
// (2, 12, 'sp12_v_b_4')
// (2, 12, 'sp4_r_v_b_5')
// (2, 13, 'neigh_op_bot_2')
// (2, 13, 'sp12_v_b_3')
// (2, 14, 'sp12_v_b_0')
// (3, 8, 'sp4_h_r_10')
// (3, 8, 'sp4_v_t_40')
// (3, 9, 'sp4_v_b_40')
// (3, 10, 'sp4_v_b_29')
// (3, 11, 'neigh_op_tnl_2')
// (3, 11, 'sp4_v_b_16')
// (3, 12, 'neigh_op_lft_2')
// (3, 12, 'sp12_h_r_15')
// (3, 12, 'sp4_v_b_5')
// (3, 13, 'neigh_op_bnl_2')
// (4, 8, 'local_g0_7')
// (4, 8, 'lutff_7/in_0')
// (4, 8, 'sp4_h_r_23')
// (4, 12, 'local_g1_0')
// (4, 12, 'lutff_7/in_0')
// (4, 12, 'sp12_h_r_16')
// (5, 8, 'sp4_h_r_34')
// (5, 12, 'sp12_h_r_19')
// (6, 8, 'sp4_h_r_47')
// (6, 12, 'sp12_h_r_20')
// (7, 8, 'sp4_h_l_47')
// (7, 12, 'sp12_h_r_23')
// (8, 12, 'sp12_h_l_23')

wire n33;
// (0, 12, 'span12_horz_9')
// (1, 12, 'local_g0_2')
// (1, 12, 'lutff_0/in_0')
// (1, 12, 'sp12_h_r_10')
// (2, 8, 'sp4_h_r_11')
// (2, 12, 'sp12_h_r_13')
// (3, 8, 'sp4_h_r_22')
// (3, 12, 'sp12_h_r_14')
// (4, 8, 'local_g3_3')
// (4, 8, 'lutff_4/in_2')
// (4, 8, 'sp4_h_r_35')
// (4, 11, 'neigh_op_tnr_5')
// (4, 12, 'neigh_op_rgt_5')
// (4, 12, 'sp12_h_r_17')
// (4, 13, 'neigh_op_bnr_5')
// (5, 8, 'sp4_h_r_46')
// (5, 9, 'sp4_r_v_b_46')
// (5, 10, 'local_g0_0')
// (5, 10, 'lutff_6/in_2')
// (5, 10, 'sp4_r_v_b_35')
// (5, 11, 'neigh_op_top_5')
// (5, 11, 'sp4_r_v_b_22')
// (5, 12, 'lutff_5/out')
// (5, 12, 'sp12_h_r_18')
// (5, 12, 'sp4_r_v_b_11')
// (5, 13, 'neigh_op_bot_5')
// (6, 8, 'sp4_h_l_46')
// (6, 8, 'sp4_v_t_46')
// (6, 9, 'sp4_v_b_46')
// (6, 10, 'sp4_v_b_35')
// (6, 11, 'neigh_op_tnl_5')
// (6, 11, 'sp4_v_b_22')
// (6, 12, 'neigh_op_lft_5')
// (6, 12, 'sp12_h_r_21')
// (6, 12, 'sp4_v_b_11')
// (6, 13, 'neigh_op_bnl_5')
// (7, 12, 'sp12_h_r_22')
// (8, 12, 'sp12_h_l_22')

reg n34 = 0;
// (0, 13, 'span12_horz_1')
// (1, 13, 'sp12_h_r_2')
// (2, 13, 'sp12_h_r_5')
// (3, 13, 'sp12_h_r_6')
// (4, 13, 'sp12_h_r_9')
// (5, 13, 'sp12_h_r_10')
// (6, 13, 'sp12_h_r_13')
// (7, 13, 'sp12_h_r_14')
// (8, 12, 'neigh_op_tnr_5')
// (8, 13, 'neigh_op_rgt_5')
// (8, 13, 'sp12_h_r_17')
// (8, 13, 'sp4_h_r_8')
// (8, 14, 'neigh_op_bnr_5')
// (9, 12, 'neigh_op_top_5')
// (9, 13, 'local_g0_5')
// (9, 13, 'lutff_5/in_2')
// (9, 13, 'lutff_5/out')
// (9, 13, 'sp12_h_r_18')
// (9, 13, 'sp4_h_r_21')
// (9, 14, 'neigh_op_bot_5')
// (10, 12, 'neigh_op_tnl_5')
// (10, 13, 'neigh_op_lft_5')
// (10, 13, 'sp12_h_r_21')
// (10, 13, 'sp4_h_r_32')
// (10, 14, 'neigh_op_bnl_5')
// (11, 10, 'sp4_r_v_b_39')
// (11, 10, 'sp4_r_v_b_45')
// (11, 11, 'local_g0_2')
// (11, 11, 'local_g1_2')
// (11, 11, 'lutff_0/in_2')
// (11, 11, 'lutff_4/in_0')
// (11, 11, 'lutff_7/in_2')
// (11, 11, 'sp4_r_v_b_26')
// (11, 11, 'sp4_r_v_b_32')
// (11, 12, 'local_g3_5')
// (11, 12, 'lutff_4/in_0')
// (11, 12, 'sp4_r_v_b_15')
// (11, 12, 'sp4_r_v_b_21')
// (11, 13, 'local_g1_6')
// (11, 13, 'lutff_1/in_2')
// (11, 13, 'sp12_h_r_22')
// (11, 13, 'sp4_h_r_45')
// (11, 13, 'sp4_r_v_b_2')
// (11, 13, 'sp4_r_v_b_8')
// (12, 9, 'sp4_v_t_39')
// (12, 9, 'sp4_v_t_45')
// (12, 10, 'sp4_v_b_39')
// (12, 10, 'sp4_v_b_45')
// (12, 11, 'sp4_v_b_26')
// (12, 11, 'sp4_v_b_32')
// (12, 12, 'sp4_v_b_15')
// (12, 12, 'sp4_v_b_21')
// (12, 13, 'sp12_h_l_22')
// (12, 13, 'sp4_h_l_45')
// (12, 13, 'sp4_v_b_2')
// (12, 13, 'sp4_v_b_8')

wire n35;
// (0, 13, 'span12_horz_2')
// (1, 12, 'neigh_op_tnr_7')
// (1, 13, 'neigh_op_rgt_7')
// (1, 13, 'sp12_h_r_5')
// (1, 13, 'sp4_h_r_2')
// (1, 14, 'neigh_op_bnr_7')
// (2, 11, 'sp4_r_v_b_39')
// (2, 12, 'neigh_op_top_7')
// (2, 12, 'sp4_r_v_b_26')
// (2, 13, 'lutff_7/out')
// (2, 13, 'sp12_h_r_6')
// (2, 13, 'sp4_h_r_15')
// (2, 13, 'sp4_r_v_b_15')
// (2, 14, 'neigh_op_bot_7')
// (2, 14, 'sp4_r_v_b_2')
// (3, 10, 'sp4_v_t_39')
// (3, 11, 'sp4_v_b_39')
// (3, 12, 'neigh_op_tnl_7')
// (3, 12, 'sp4_v_b_26')
// (3, 13, 'neigh_op_lft_7')
// (3, 13, 'sp12_h_r_9')
// (3, 13, 'sp4_h_r_26')
// (3, 13, 'sp4_v_b_15')
// (3, 14, 'neigh_op_bnl_7')
// (3, 14, 'sp4_h_r_2')
// (3, 14, 'sp4_v_b_2')
// (4, 10, 'sp4_r_v_b_45')
// (4, 11, 'sp4_r_v_b_32')
// (4, 12, 'sp4_r_v_b_21')
// (4, 13, 'sp12_h_r_10')
// (4, 13, 'sp4_h_r_39')
// (4, 13, 'sp4_r_v_b_8')
// (4, 14, 'local_g0_7')
// (4, 14, 'lutff_5/in_2')
// (4, 14, 'sp4_h_r_15')
// (5, 9, 'sp4_h_r_1')
// (5, 9, 'sp4_v_t_45')
// (5, 10, 'sp4_v_b_45')
// (5, 11, 'sp4_v_b_32')
// (5, 12, 'local_g0_5')
// (5, 12, 'lutff_5/in_0')
// (5, 12, 'sp4_v_b_21')
// (5, 13, 'sp12_h_r_13')
// (5, 13, 'sp4_h_l_39')
// (5, 13, 'sp4_v_b_8')
// (5, 14, 'sp4_h_r_26')
// (6, 9, 'sp4_h_r_12')
// (6, 11, 'sp4_r_v_b_45')
// (6, 12, 'local_g0_3')
// (6, 12, 'lutff_3/in_0')
// (6, 12, 'sp4_r_v_b_32')
// (6, 13, 'sp12_h_r_14')
// (6, 13, 'sp4_r_v_b_21')
// (6, 14, 'sp4_h_r_39')
// (6, 14, 'sp4_r_v_b_8')
// (7, 9, 'sp4_h_r_25')
// (7, 10, 'sp4_v_t_45')
// (7, 11, 'sp4_v_b_45')
// (7, 12, 'local_g2_0')
// (7, 12, 'local_g3_0')
// (7, 12, 'lutff_2/in_3')
// (7, 12, 'lutff_3/in_3')
// (7, 12, 'lutff_6/in_3')
// (7, 12, 'sp4_v_b_32')
// (7, 13, 'sp12_h_r_17')
// (7, 13, 'sp4_v_b_21')
// (7, 14, 'sp4_h_l_39')
// (7, 14, 'sp4_v_b_8')
// (8, 9, 'sp4_h_r_36')
// (8, 10, 'sp4_r_v_b_36')
// (8, 11, 'sp4_r_v_b_25')
// (8, 12, 'local_g2_4')
// (8, 12, 'lutff_0/in_0')
// (8, 12, 'sp4_r_v_b_12')
// (8, 13, 'local_g1_2')
// (8, 13, 'lutff_2/in_3')
// (8, 13, 'lutff_4/in_3')
// (8, 13, 'sp12_h_r_18')
// (8, 13, 'sp4_r_v_b_1')
// (9, 9, 'sp4_h_l_36')
// (9, 9, 'sp4_v_t_36')
// (9, 10, 'sp4_v_b_36')
// (9, 11, 'sp4_v_b_25')
// (9, 12, 'sp4_v_b_12')
// (9, 13, 'sp12_h_r_21')
// (9, 13, 'sp4_v_b_1')
// (10, 13, 'sp12_h_r_22')
// (11, 13, 'sp12_h_l_22')

wire n36;
// (0, 14, 'span12_horz_0')
// (1, 14, 'sp12_h_r_3')
// (2, 14, 'sp12_h_r_4')
// (3, 14, 'sp12_h_r_7')
// (4, 14, 'sp12_h_r_8')
// (5, 13, 'neigh_op_tnr_2')
// (5, 14, 'neigh_op_rgt_2')
// (5, 14, 'sp12_h_r_11')
// (5, 15, 'neigh_op_bnr_2')
// (6, 13, 'neigh_op_top_2')
// (6, 14, 'local_g0_2')
// (6, 14, 'lutff_2/out')
// (6, 14, 'lutff_5/in_1')
// (6, 14, 'lutff_7/in_1')
// (6, 14, 'sp12_h_r_12')
// (6, 15, 'neigh_op_bot_2')
// (7, 13, 'neigh_op_tnl_2')
// (7, 14, 'neigh_op_lft_2')
// (7, 14, 'sp12_h_r_15')
// (7, 14, 'sp4_h_r_9')
// (7, 15, 'neigh_op_bnl_2')
// (8, 14, 'local_g0_4')
// (8, 14, 'local_g1_0')
// (8, 14, 'lutff_3/in_2')
// (8, 14, 'lutff_4/in_3')
// (8, 14, 'lutff_7/in_3')
// (8, 14, 'sp12_h_r_16')
// (8, 14, 'sp4_h_r_20')
// (9, 14, 'sp12_h_r_19')
// (9, 14, 'sp4_h_r_33')
// (10, 14, 'sp12_h_r_20')
// (10, 14, 'sp4_h_r_44')
// (11, 14, 'sp12_h_r_23')
// (11, 14, 'sp4_h_l_44')
// (12, 14, 'sp12_h_l_23')

wire rst;
// (0, 14, 'span4_horz_31')
// (0, 14, 'span4_horz_7')
// (1, 11, 'sp4_r_v_b_47')
// (1, 12, 'sp4_r_v_b_34')
// (1, 13, 'sp4_r_v_b_23')
// (1, 14, 'sp4_h_r_18')
// (1, 14, 'sp4_h_r_42')
// (1, 14, 'sp4_r_v_b_10')
// (2, 10, 'sp4_v_t_47')
// (2, 11, 'sp4_v_b_47')
// (2, 12, 'sp12_h_r_0')
// (2, 12, 'sp12_v_t_23')
// (2, 12, 'sp4_v_b_34')
// (2, 13, 'sp12_v_b_23')
// (2, 13, 'sp4_v_b_23')
// (2, 14, 'sp12_v_b_20')
// (2, 14, 'sp4_h_l_42')
// (2, 14, 'sp4_h_r_31')
// (2, 14, 'sp4_h_r_4')
// (2, 14, 'sp4_v_b_10')
// (2, 15, 'local_g2_3')
// (2, 15, 'lutff_2/in_3')
// (2, 15, 'lutff_6/in_3')
// (2, 15, 'sp12_v_b_19')
// (2, 16, 'sp12_v_b_16')
// (2, 17, 'span12_vert_15')
// (3, 11, 'sp4_r_v_b_42')
// (3, 12, 'sp12_h_r_3')
// (3, 12, 'sp4_r_v_b_31')
// (3, 13, 'sp4_r_v_b_18')
// (3, 14, 'sp4_h_r_17')
// (3, 14, 'sp4_h_r_42')
// (3, 14, 'sp4_r_v_b_7')
// (4, 10, 'sp4_v_t_42')
// (4, 11, 'sp4_v_b_42')
// (4, 12, 'sp12_h_r_4')
// (4, 12, 'sp4_v_b_31')
// (4, 13, 'local_g0_2')
// (4, 13, 'lutff_7/in_1')
// (4, 13, 'sp4_v_b_18')
// (4, 14, 'local_g2_4')
// (4, 14, 'lutff_global/s_r')
// (4, 14, 'sp4_h_l_42')
// (4, 14, 'sp4_h_r_28')
// (4, 14, 'sp4_v_b_7')
// (5, 12, 'sp12_h_r_7')
// (5, 14, 'sp4_h_r_41')
// (5, 15, 'local_g3_1')
// (5, 15, 'local_g3_4')
// (5, 15, 'lutff_0/in_1')
// (5, 15, 'lutff_2/in_3')
// (5, 15, 'lutff_7/in_3')
// (5, 15, 'sp4_r_v_b_41')
// (5, 15, 'sp4_r_v_b_44')
// (5, 16, 'sp4_r_v_b_28')
// (5, 16, 'sp4_r_v_b_33')
// (6, 12, 'sp12_h_r_8')
// (6, 14, 'sp4_h_l_41')
// (6, 14, 'sp4_v_t_41')
// (6, 14, 'sp4_v_t_44')
// (6, 15, 'sp4_v_b_41')
// (6, 15, 'sp4_v_b_44')
// (6, 16, 'sp4_v_b_28')
// (6, 16, 'sp4_v_b_33')
// (6, 17, 'span4_vert_17')
// (6, 17, 'span4_vert_20')
// (7, 12, 'sp12_h_r_11')
// (8, 12, 'sp12_h_r_12')
// (9, 12, 'sp12_h_r_15')
// (9, 13, 'sp4_r_v_b_41')
// (9, 14, 'local_g0_4')
// (9, 14, 'lutff_1/in_3')
// (9, 14, 'sp4_r_v_b_28')
// (9, 15, 'sp4_r_v_b_17')
// (9, 16, 'sp4_r_v_b_4')
// (10, 12, 'sp12_h_r_16')
// (10, 12, 'sp4_h_r_4')
// (10, 12, 'sp4_v_t_41')
// (10, 13, 'sp4_v_b_41')
// (10, 14, 'sp4_v_b_28')
// (10, 15, 'sp4_v_b_17')
// (10, 16, 'sp4_v_b_4')
// (11, 12, 'local_g1_1')
// (11, 12, 'lutff_3/in_3')
// (11, 12, 'lutff_5/in_3')
// (11, 12, 'sp12_h_r_19')
// (11, 12, 'sp4_h_r_17')
// (12, 11, 'neigh_op_tnr_2')
// (12, 11, 'neigh_op_tnr_6')
// (12, 12, 'local_g3_2')
// (12, 12, 'lutff_0/in_3')
// (12, 12, 'neigh_op_rgt_2')
// (12, 12, 'neigh_op_rgt_6')
// (12, 12, 'sp12_h_r_20')
// (12, 12, 'sp4_h_r_28')
// (12, 13, 'neigh_op_bnr_2')
// (12, 13, 'neigh_op_bnr_6')
// (13, 12, 'io_1/D_IN_0')
// (13, 12, 'io_1/PAD')
// (13, 12, 'span12_horz_20')
// (13, 12, 'span4_horz_28')

reg n38 = 0;
// (0, 15, 'span12_horz_0')
// (0, 15, 'span12_horz_16')
// (1, 14, 'neigh_op_tnr_6')
// (1, 15, 'neigh_op_rgt_6')
// (1, 15, 'sp12_h_r_19')
// (1, 15, 'sp12_h_r_3')
// (1, 16, 'neigh_op_bnr_6')
// (2, 9, 'sp12_v_t_23')
// (2, 10, 'sp12_v_b_23')
// (2, 11, 'local_g2_4')
// (2, 11, 'lutff_2/in_2')
// (2, 11, 'sp12_v_b_20')
// (2, 12, 'local_g2_3')
// (2, 12, 'lutff_1/in_2')
// (2, 12, 'sp12_v_b_19')
// (2, 13, 'local_g2_0')
// (2, 13, 'lutff_7/in_3')
// (2, 13, 'sp12_v_b_16')
// (2, 13, 'sp4_r_v_b_37')
// (2, 14, 'neigh_op_top_6')
// (2, 14, 'sp12_v_b_15')
// (2, 14, 'sp4_r_v_b_24')
// (2, 15, 'local_g1_6')
// (2, 15, 'lutff_2/in_1')
// (2, 15, 'lutff_6/in_1')
// (2, 15, 'lutff_6/out')
// (2, 15, 'sp12_h_r_20')
// (2, 15, 'sp12_h_r_4')
// (2, 15, 'sp12_v_b_12')
// (2, 15, 'sp4_r_v_b_13')
// (2, 16, 'neigh_op_bot_6')
// (2, 16, 'sp12_v_b_11')
// (2, 16, 'sp4_r_v_b_0')
// (2, 17, 'span12_vert_8')
// (3, 12, 'sp4_h_r_0')
// (3, 12, 'sp4_r_v_b_37')
// (3, 12, 'sp4_v_t_37')
// (3, 13, 'sp4_r_v_b_24')
// (3, 13, 'sp4_v_b_37')
// (3, 14, 'neigh_op_tnl_6')
// (3, 14, 'sp4_r_v_b_13')
// (3, 14, 'sp4_v_b_24')
// (3, 15, 'neigh_op_lft_6')
// (3, 15, 'sp12_h_r_23')
// (3, 15, 'sp12_h_r_7')
// (3, 15, 'sp4_r_v_b_0')
// (3, 15, 'sp4_v_b_13')
// (3, 16, 'neigh_op_bnl_6')
// (3, 16, 'sp4_v_b_0')
// (4, 3, 'sp12_v_t_23')
// (4, 4, 'sp12_v_b_23')
// (4, 5, 'sp12_v_b_20')
// (4, 6, 'sp12_v_b_19')
// (4, 7, 'sp12_v_b_16')
// (4, 8, 'sp12_v_b_15')
// (4, 9, 'sp12_v_b_12')
// (4, 10, 'sp12_v_b_11')
// (4, 11, 'local_g3_0')
// (4, 11, 'lutff_2/in_3')
// (4, 11, 'sp12_v_b_8')
// (4, 11, 'sp4_h_r_5')
// (4, 11, 'sp4_v_t_37')
// (4, 12, 'local_g2_7')
// (4, 12, 'local_g3_7')
// (4, 12, 'lutff_1/in_2')
// (4, 12, 'lutff_2/in_2')
// (4, 12, 'lutff_3/in_2')
// (4, 12, 'sp12_v_b_7')
// (4, 12, 'sp4_h_r_13')
// (4, 12, 'sp4_r_v_b_37')
// (4, 12, 'sp4_v_b_37')
// (4, 13, 'sp12_v_b_4')
// (4, 13, 'sp4_r_v_b_24')
// (4, 13, 'sp4_v_b_24')
// (4, 14, 'sp12_v_b_3')
// (4, 14, 'sp4_r_v_b_13')
// (4, 14, 'sp4_v_b_13')
// (4, 15, 'local_g1_0')
// (4, 15, 'lutff_0/in_3')
// (4, 15, 'sp12_h_l_23')
// (4, 15, 'sp12_h_r_8')
// (4, 15, 'sp12_v_b_0')
// (4, 15, 'sp4_r_v_b_0')
// (4, 15, 'sp4_v_b_0')
// (5, 11, 'local_g0_0')
// (5, 11, 'local_g1_0')
// (5, 11, 'lutff_0/in_2')
// (5, 11, 'lutff_1/in_2')
// (5, 11, 'lutff_3/in_2')
// (5, 11, 'lutff_4/in_2')
// (5, 11, 'sp4_h_r_16')
// (5, 11, 'sp4_v_t_37')
// (5, 12, 'local_g2_0')
// (5, 12, 'local_g3_0')
// (5, 12, 'lutff_0/in_2')
// (5, 12, 'lutff_1/in_2')
// (5, 12, 'sp4_h_r_24')
// (5, 12, 'sp4_v_b_37')
// (5, 13, 'sp4_v_b_24')
// (5, 14, 'local_g0_5')
// (5, 14, 'lutff_7/in_2')
// (5, 14, 'sp4_v_b_13')
// (5, 15, 'sp12_h_r_11')
// (5, 15, 'sp4_h_r_7')
// (5, 15, 'sp4_v_b_0')
// (6, 11, 'local_g2_5')
// (6, 11, 'local_g3_5')
// (6, 11, 'lutff_1/in_2')
// (6, 11, 'lutff_3/in_2')
// (6, 11, 'lutff_6/in_2')
// (6, 11, 'sp4_h_r_29')
// (6, 12, 'sp4_h_r_37')
// (6, 15, 'sp12_h_r_12')
// (6, 15, 'sp4_h_r_18')
// (7, 11, 'sp4_h_r_40')
// (7, 12, 'sp4_h_l_37')
// (7, 15, 'sp12_h_r_15')
// (7, 15, 'sp4_h_r_31')
// (8, 11, 'sp4_h_l_40')
// (8, 15, 'sp12_h_r_16')
// (8, 15, 'sp4_h_r_42')
// (9, 15, 'sp12_h_r_19')
// (9, 15, 'sp4_h_l_42')
// (10, 15, 'sp12_h_r_20')
// (11, 15, 'sp12_h_r_23')
// (12, 15, 'sp12_h_l_23')

wire n39;
// (0, 15, 'span12_horz_2')
// (1, 15, 'sp12_h_r_5')
// (2, 15, 'sp12_h_r_6')
// (3, 14, 'neigh_op_tnr_1')
// (3, 15, 'neigh_op_rgt_1')
// (3, 15, 'sp12_h_r_9')
// (3, 16, 'neigh_op_bnr_1')
// (4, 14, 'neigh_op_top_1')
// (4, 15, 'local_g2_1')
// (4, 15, 'local_g3_1')
// (4, 15, 'lutff_1/out')
// (4, 15, 'lutff_3/in_1')
// (4, 15, 'lutff_7/in_0')
// (4, 15, 'sp12_h_r_10')
// (4, 16, 'neigh_op_bot_1')
// (5, 14, 'neigh_op_tnl_1')
// (5, 15, 'neigh_op_lft_1')
// (5, 15, 'sp12_h_r_13')
// (5, 16, 'neigh_op_bnl_1')
// (6, 15, 'sp12_h_r_14')
// (7, 15, 'sp12_h_r_17')
// (8, 12, 'sp4_r_v_b_38')
// (8, 13, 'sp4_r_v_b_27')
// (8, 14, 'sp4_r_v_b_14')
// (8, 15, 'sp12_h_r_18')
// (8, 15, 'sp4_r_v_b_3')
// (9, 11, 'sp4_v_t_38')
// (9, 12, 'sp4_v_b_38')
// (9, 13, 'sp4_v_b_27')
// (9, 14, 'local_g0_6')
// (9, 14, 'lutff_1/in_1')
// (9, 14, 'sp4_v_b_14')
// (9, 15, 'sp12_h_r_21')
// (9, 15, 'sp4_h_r_10')
// (9, 15, 'sp4_v_b_3')
// (10, 15, 'sp12_h_r_22')
// (10, 15, 'sp4_h_r_23')
// (11, 3, 'sp12_v_t_22')
// (11, 4, 'sp12_v_b_22')
// (11, 5, 'sp12_v_b_21')
// (11, 6, 'sp12_v_b_18')
// (11, 7, 'sp12_v_b_17')
// (11, 8, 'sp12_v_b_14')
// (11, 9, 'sp12_v_b_13')
// (11, 10, 'sp12_v_b_10')
// (11, 11, 'sp12_v_b_9')
// (11, 12, 'local_g2_6')
// (11, 12, 'lutff_5/in_1')
// (11, 12, 'sp12_v_b_6')
// (11, 13, 'sp12_v_b_5')
// (11, 14, 'sp12_v_b_2')
// (11, 15, 'sp12_h_l_22')
// (11, 15, 'sp12_v_b_1')
// (11, 15, 'sp4_h_r_34')
// (12, 15, 'sp4_h_r_47')
// (13, 15, 'span4_horz_47')

reg n40 = 0;
// (1, 2, 'neigh_op_tnr_3')
// (1, 3, 'neigh_op_rgt_3')
// (1, 4, 'neigh_op_bnr_3')
// (2, 2, 'neigh_op_top_3')
// (2, 3, 'lutff_3/out')
// (2, 3, 'sp4_h_r_6')
// (2, 4, 'neigh_op_bot_3')
// (3, 2, 'neigh_op_tnl_3')
// (3, 3, 'neigh_op_lft_3')
// (3, 3, 'sp4_h_r_19')
// (3, 4, 'neigh_op_bnl_3')
// (4, 3, 'sp4_h_r_30')
// (5, 3, 'local_g2_3')
// (5, 3, 'lutff_1/in_0')
// (5, 3, 'sp4_h_r_43')
// (6, 3, 'sp4_h_l_43')

reg n41 = 0;
// (1, 3, 'neigh_op_tnr_0')
// (1, 4, 'neigh_op_rgt_0')
// (1, 5, 'neigh_op_bnr_0')
// (2, 3, 'neigh_op_top_0')
// (2, 4, 'lutff_0/out')
// (2, 5, 'local_g0_0')
// (2, 5, 'lutff_2/in_0')
// (2, 5, 'neigh_op_bot_0')
// (3, 3, 'neigh_op_tnl_0')
// (3, 4, 'neigh_op_lft_0')
// (3, 5, 'neigh_op_bnl_0')

reg n42 = 0;
// (1, 3, 'sp4_r_v_b_42')
// (1, 4, 'sp4_r_v_b_31')
// (1, 5, 'sp4_r_v_b_18')
// (1, 6, 'sp4_r_v_b_7')
// (2, 0, 'span12_vert_21')
// (2, 1, 'sp12_v_b_21')
// (2, 2, 'sp12_v_b_18')
// (2, 2, 'sp4_v_t_42')
// (2, 3, 'sp12_v_b_17')
// (2, 3, 'sp4_v_b_42')
// (2, 4, 'sp12_v_b_14')
// (2, 4, 'sp4_v_b_31')
// (2, 5, 'sp12_v_b_13')
// (2, 5, 'sp4_v_b_18')
// (2, 6, 'sp12_v_b_10')
// (2, 6, 'sp4_h_r_7')
// (2, 6, 'sp4_v_b_7')
// (2, 7, 'local_g2_1')
// (2, 7, 'local_g3_1')
// (2, 7, 'lutff_0/in_3')
// (2, 7, 'lutff_7/in_3')
// (2, 7, 'sp12_v_b_9')
// (2, 8, 'local_g3_6')
// (2, 8, 'lutff_5/in_2')
// (2, 8, 'sp12_v_b_6')
// (2, 9, 'sp12_v_b_5')
// (2, 10, 'sp12_v_b_2')
// (2, 11, 'sp12_h_r_1')
// (2, 11, 'sp12_v_b_1')
// (3, 6, 'sp4_h_r_18')
// (3, 11, 'sp12_h_r_2')
// (4, 6, 'sp4_h_r_31')
// (4, 11, 'sp12_h_r_5')
// (5, 3, 'sp4_r_v_b_42')
// (5, 4, 'sp4_r_v_b_31')
// (5, 5, 'sp4_r_v_b_18')
// (5, 6, 'local_g2_2')
// (5, 6, 'lutff_0/in_2')
// (5, 6, 'lutff_3/in_3')
// (5, 6, 'lutff_7/in_3')
// (5, 6, 'sp4_h_r_42')
// (5, 6, 'sp4_r_v_b_7')
// (5, 7, 'local_g2_6')
// (5, 7, 'lutff_0/in_2')
// (5, 7, 'sp4_r_v_b_37')
// (5, 7, 'sp4_r_v_b_38')
// (5, 7, 'sp4_r_v_b_47')
// (5, 8, 'sp4_r_v_b_24')
// (5, 8, 'sp4_r_v_b_27')
// (5, 8, 'sp4_r_v_b_34')
// (5, 9, 'local_g2_5')
// (5, 9, 'local_g2_6')
// (5, 9, 'lutff_1/in_2')
// (5, 9, 'lutff_5/in_3')
// (5, 9, 'lutff_6/in_3')
// (5, 9, 'sp4_r_v_b_13')
// (5, 9, 'sp4_r_v_b_14')
// (5, 9, 'sp4_r_v_b_23')
// (5, 10, 'sp4_r_v_b_0')
// (5, 10, 'sp4_r_v_b_10')
// (5, 10, 'sp4_r_v_b_3')
// (5, 11, 'sp12_h_r_6')
// (6, 2, 'sp4_v_t_42')
// (6, 3, 'local_g2_2')
// (6, 3, 'local_g3_2')
// (6, 3, 'lutff_0/in_2')
// (6, 3, 'lutff_1/in_3')
// (6, 3, 'lutff_2/in_3')
// (6, 3, 'sp4_v_b_42')
// (6, 4, 'sp4_v_b_31')
// (6, 5, 'sp4_v_b_18')
// (6, 6, 'local_g0_7')
// (6, 6, 'lutff_1/in_2')
// (6, 6, 'sp4_h_l_42')
// (6, 6, 'sp4_v_b_7')
// (6, 6, 'sp4_v_t_37')
// (6, 6, 'sp4_v_t_38')
// (6, 6, 'sp4_v_t_47')
// (6, 7, 'sp4_v_b_37')
// (6, 7, 'sp4_v_b_38')
// (6, 7, 'sp4_v_b_47')
// (6, 8, 'local_g2_0')
// (6, 8, 'local_g3_0')
// (6, 8, 'lutff_3/in_3')
// (6, 8, 'lutff_6/in_3')
// (6, 8, 'sp4_v_b_24')
// (6, 8, 'sp4_v_b_27')
// (6, 8, 'sp4_v_b_34')
// (6, 9, 'local_g0_6')
// (6, 9, 'local_g0_7')
// (6, 9, 'lutff_0/in_3')
// (6, 9, 'lutff_1/in_3')
// (6, 9, 'sp4_v_b_13')
// (6, 9, 'sp4_v_b_14')
// (6, 9, 'sp4_v_b_23')
// (6, 10, 'sp4_v_b_0')
// (6, 10, 'sp4_v_b_10')
// (6, 10, 'sp4_v_b_3')
// (6, 11, 'sp12_h_r_9')
// (7, 1, 'local_g0_3')
// (7, 1, 'lutff_6/in_3')
// (7, 1, 'sp4_h_r_11')
// (7, 11, 'sp12_h_r_10')
// (8, 1, 'sp4_h_r_22')
// (8, 7, 'local_g1_3')
// (8, 7, 'lutff_0/in_2')
// (8, 7, 'sp4_h_r_11')
// (8, 11, 'sp12_h_r_13')
// (9, 1, 'sp4_h_r_35')
// (9, 7, 'sp4_h_r_22')
// (9, 11, 'sp12_h_r_14')
// (10, 1, 'sp4_h_r_46')
// (10, 2, 'sp4_r_v_b_40')
// (10, 3, 'sp4_r_v_b_29')
// (10, 4, 'sp4_r_v_b_16')
// (10, 5, 'sp4_r_v_b_5')
// (10, 6, 'sp4_r_v_b_44')
// (10, 7, 'sp4_h_r_35')
// (10, 7, 'sp4_r_v_b_33')
// (10, 8, 'sp4_r_v_b_20')
// (10, 9, 'sp4_r_v_b_9')
// (10, 10, 'neigh_op_tnr_5')
// (10, 11, 'neigh_op_rgt_5')
// (10, 11, 'sp12_h_r_17')
// (10, 12, 'neigh_op_bnr_5')
// (11, 1, 'sp4_h_l_46')
// (11, 1, 'sp4_v_t_40')
// (11, 2, 'sp4_v_b_40')
// (11, 3, 'sp4_v_b_29')
// (11, 4, 'sp12_v_t_22')
// (11, 4, 'sp4_v_b_16')
// (11, 5, 'sp12_v_b_22')
// (11, 5, 'sp4_v_b_5')
// (11, 5, 'sp4_v_t_44')
// (11, 6, 'sp12_v_b_21')
// (11, 6, 'sp4_v_b_44')
// (11, 7, 'local_g3_1')
// (11, 7, 'local_g3_2')
// (11, 7, 'lutff_0/in_3')
// (11, 7, 'lutff_7/in_3')
// (11, 7, 'sp12_v_b_18')
// (11, 7, 'sp4_h_r_46')
// (11, 7, 'sp4_v_b_33')
// (11, 8, 'sp12_v_b_17')
// (11, 8, 'sp4_r_v_b_46')
// (11, 8, 'sp4_v_b_20')
// (11, 9, 'local_g1_1')
// (11, 9, 'local_g3_6')
// (11, 9, 'lutff_0/in_2')
// (11, 9, 'lutff_1/in_3')
// (11, 9, 'lutff_2/in_3')
// (11, 9, 'sp12_v_b_14')
// (11, 9, 'sp4_r_v_b_35')
// (11, 9, 'sp4_v_b_9')
// (11, 10, 'neigh_op_top_5')
// (11, 10, 'sp12_v_b_13')
// (11, 10, 'sp4_r_v_b_22')
// (11, 11, 'lutff_5/out')
// (11, 11, 'sp12_h_r_18')
// (11, 11, 'sp12_v_b_10')
// (11, 11, 'sp4_r_v_b_11')
// (11, 12, 'neigh_op_bot_5')
// (11, 12, 'sp12_v_b_9')
// (11, 13, 'sp12_v_b_6')
// (11, 14, 'sp12_v_b_5')
// (11, 15, 'sp12_v_b_2')
// (11, 16, 'sp12_v_b_1')
// (12, 7, 'sp4_h_l_46')
// (12, 7, 'sp4_v_t_46')
// (12, 8, 'sp4_v_b_46')
// (12, 9, 'sp4_v_b_35')
// (12, 10, 'neigh_op_tnl_5')
// (12, 10, 'sp4_v_b_22')
// (12, 11, 'neigh_op_lft_5')
// (12, 11, 'sp12_h_r_21')
// (12, 11, 'sp4_v_b_11')
// (12, 12, 'neigh_op_bnl_5')
// (13, 11, 'span12_horz_21')

reg n43 = 0;
// (1, 4, 'neigh_op_tnr_1')
// (1, 5, 'neigh_op_rgt_1')
// (1, 6, 'neigh_op_bnr_1')
// (2, 2, 'sp4_r_v_b_38')
// (2, 3, 'local_g0_3')
// (2, 3, 'lutff_3/in_0')
// (2, 3, 'sp4_r_v_b_27')
// (2, 4, 'neigh_op_top_1')
// (2, 4, 'sp4_r_v_b_14')
// (2, 5, 'lutff_1/out')
// (2, 5, 'sp4_r_v_b_3')
// (2, 6, 'neigh_op_bot_1')
// (3, 1, 'sp4_v_t_38')
// (3, 2, 'sp4_v_b_38')
// (3, 3, 'sp4_v_b_27')
// (3, 4, 'neigh_op_tnl_1')
// (3, 4, 'sp4_v_b_14')
// (3, 5, 'neigh_op_lft_1')
// (3, 5, 'sp4_v_b_3')
// (3, 6, 'neigh_op_bnl_1')

reg n44 = 0;
// (1, 4, 'neigh_op_tnr_2')
// (1, 5, 'neigh_op_rgt_2')
// (1, 5, 'sp4_h_r_9')
// (1, 6, 'neigh_op_bnr_2')
// (2, 4, 'neigh_op_top_2')
// (2, 5, 'lutff_2/out')
// (2, 5, 'sp4_h_r_20')
// (2, 6, 'neigh_op_bot_2')
// (3, 4, 'neigh_op_tnl_2')
// (3, 5, 'neigh_op_lft_2')
// (3, 5, 'sp4_h_r_33')
// (3, 6, 'neigh_op_bnl_2')
// (4, 5, 'sp4_h_r_44')
// (4, 6, 'sp4_r_v_b_44')
// (4, 7, 'local_g2_1')
// (4, 7, 'lutff_1/in_0')
// (4, 7, 'sp4_r_v_b_33')
// (4, 8, 'sp4_r_v_b_20')
// (4, 9, 'sp4_r_v_b_9')
// (4, 10, 'sp4_r_v_b_38')
// (4, 11, 'sp4_r_v_b_27')
// (4, 12, 'local_g2_6')
// (4, 12, 'lutff_1/in_3')
// (4, 12, 'sp4_r_v_b_14')
// (4, 13, 'sp4_r_v_b_3')
// (5, 5, 'sp4_h_l_44')
// (5, 5, 'sp4_v_t_44')
// (5, 6, 'sp4_v_b_44')
// (5, 7, 'sp4_v_b_33')
// (5, 8, 'sp4_v_b_20')
// (5, 9, 'sp4_h_r_3')
// (5, 9, 'sp4_v_b_9')
// (5, 9, 'sp4_v_t_38')
// (5, 10, 'sp4_v_b_38')
// (5, 11, 'sp4_v_b_27')
// (5, 12, 'sp4_v_b_14')
// (5, 13, 'sp4_v_b_3')
// (6, 9, 'sp4_h_r_14')
// (7, 9, 'sp4_h_r_27')
// (8, 9, 'sp4_h_r_38')
// (9, 9, 'sp4_h_l_38')

reg n45 = 0;
// (1, 6, 'neigh_op_tnr_0')
// (1, 7, 'neigh_op_rgt_0')
// (1, 8, 'neigh_op_bnr_0')
// (2, 6, 'neigh_op_top_0')
// (2, 7, 'local_g2_0')
// (2, 7, 'lutff_0/out')
// (2, 7, 'lutff_7/in_1')
// (2, 8, 'neigh_op_bot_0')
// (3, 6, 'neigh_op_tnl_0')
// (3, 7, 'neigh_op_lft_0')
// (3, 8, 'neigh_op_bnl_0')

reg n46 = 0;
// (1, 6, 'neigh_op_tnr_7')
// (1, 7, 'neigh_op_rgt_7')
// (1, 7, 'sp4_h_r_3')
// (1, 8, 'neigh_op_bnr_7')
// (2, 6, 'neigh_op_top_7')
// (2, 7, 'lutff_7/out')
// (2, 7, 'sp4_h_r_14')
// (2, 8, 'neigh_op_bot_7')
// (3, 6, 'neigh_op_tnl_7')
// (3, 7, 'neigh_op_lft_7')
// (3, 7, 'sp4_h_r_27')
// (3, 8, 'neigh_op_bnl_7')
// (4, 4, 'sp4_r_v_b_44')
// (4, 5, 'sp4_r_v_b_33')
// (4, 6, 'sp4_r_v_b_20')
// (4, 7, 'sp4_h_r_38')
// (4, 7, 'sp4_r_v_b_9')
// (5, 3, 'sp4_v_t_44')
// (5, 4, 'sp4_v_b_44')
// (5, 5, 'sp4_v_b_33')
// (5, 6, 'sp4_v_b_20')
// (5, 7, 'local_g0_1')
// (5, 7, 'lutff_0/in_1')
// (5, 7, 'sp4_h_l_38')
// (5, 7, 'sp4_v_b_9')

wire n47;
// (1, 6, 'sp12_h_r_0')
// (2, 6, 'sp12_h_r_3')
// (3, 6, 'sp12_h_r_4')
// (4, 5, 'neigh_op_tnr_0')
// (4, 6, 'neigh_op_rgt_0')
// (4, 6, 'sp12_h_r_7')
// (4, 7, 'neigh_op_bnr_0')
// (5, 5, 'neigh_op_top_0')
// (5, 6, 'lutff_0/out')
// (5, 6, 'sp12_h_r_8')
// (5, 7, 'neigh_op_bot_0')
// (6, 5, 'neigh_op_tnl_0')
// (6, 6, 'neigh_op_lft_0')
// (6, 6, 'sp12_h_r_11')
// (6, 7, 'neigh_op_bnl_0')
// (7, 6, 'sp12_h_r_12')
// (8, 6, 'local_g0_7')
// (8, 6, 'local_g1_7')
// (8, 6, 'lutff_2/in_0')
// (8, 6, 'lutff_4/in_1')
// (8, 6, 'sp12_h_r_15')
// (9, 6, 'sp12_h_r_16')
// (10, 6, 'sp12_h_r_19')
// (11, 6, 'sp12_h_r_20')
// (12, 6, 'sp12_h_r_23')
// (13, 6, 'span12_horz_23')

wire n48;
// (1, 7, 'neigh_op_tnr_5')
// (1, 8, 'neigh_op_rgt_5')
// (1, 9, 'neigh_op_bnr_5')
// (2, 7, 'neigh_op_top_5')
// (2, 8, 'lutff_5/out')
// (2, 8, 'sp4_h_r_10')
// (2, 9, 'neigh_op_bot_5')
// (3, 7, 'neigh_op_tnl_5')
// (3, 8, 'neigh_op_lft_5')
// (3, 8, 'sp4_h_r_23')
// (3, 9, 'neigh_op_bnl_5')
// (4, 8, 'sp4_h_r_34')
// (5, 5, 'sp4_r_v_b_47')
// (5, 6, 'sp4_r_v_b_34')
// (5, 7, 'sp4_r_v_b_23')
// (5, 8, 'sp4_h_r_47')
// (5, 8, 'sp4_r_v_b_10')
// (6, 4, 'sp4_v_t_47')
// (6, 5, 'sp4_v_b_47')
// (6, 6, 'sp4_v_b_34')
// (6, 7, 'local_g0_7')
// (6, 7, 'local_g1_7')
// (6, 7, 'lutff_0/in_0')
// (6, 7, 'lutff_4/in_1')
// (6, 7, 'sp4_v_b_23')
// (6, 8, 'sp4_h_l_47')
// (6, 8, 'sp4_v_b_10')

reg n49 = 0;
// (1, 7, 'neigh_op_tnr_6')
// (1, 8, 'neigh_op_rgt_6')
// (1, 9, 'neigh_op_bnr_6')
// (2, 7, 'local_g1_6')
// (2, 7, 'lutff_0/in_1')
// (2, 7, 'neigh_op_top_6')
// (2, 8, 'lutff_6/out')
// (2, 9, 'neigh_op_bot_6')
// (3, 7, 'neigh_op_tnl_6')
// (3, 8, 'neigh_op_lft_6')
// (3, 9, 'neigh_op_bnl_6')

reg n50 = 0;
// (1, 7, 'sp12_h_r_1')
// (2, 7, 'sp12_h_r_2')
// (3, 7, 'sp12_h_r_5')
// (4, 7, 'sp12_h_r_6')
// (5, 7, 'sp12_h_r_9')
// (6, 7, 'sp12_h_r_10')
// (7, 6, 'neigh_op_tnr_3')
// (7, 7, 'neigh_op_rgt_3')
// (7, 7, 'sp12_h_r_13')
// (7, 8, 'neigh_op_bnr_3')
// (8, 6, 'neigh_op_top_3')
// (8, 7, 'local_g0_3')
// (8, 7, 'lutff_2/in_1')
// (8, 7, 'lutff_3/out')
// (8, 7, 'sp12_h_r_14')
// (8, 8, 'neigh_op_bot_3')
// (9, 6, 'neigh_op_tnl_3')
// (9, 7, 'neigh_op_lft_3')
// (9, 7, 'sp12_h_r_17')
// (9, 8, 'neigh_op_bnl_3')
// (10, 7, 'sp12_h_r_18')
// (11, 7, 'local_g0_5')
// (11, 7, 'lutff_7/in_2')
// (11, 7, 'sp12_h_r_21')
// (12, 7, 'sp12_h_r_22')
// (13, 7, 'span12_horz_22')

reg n51 = 0;
// (1, 7, 'sp4_h_r_7')
// (2, 7, 'sp4_h_r_18')
// (3, 6, 'neigh_op_tnr_5')
// (3, 7, 'neigh_op_rgt_5')
// (3, 7, 'sp4_h_r_31')
// (3, 8, 'neigh_op_bnr_5')
// (4, 6, 'neigh_op_top_5')
// (4, 7, 'lutff_5/out')
// (4, 7, 'sp4_h_r_42')
// (4, 8, 'neigh_op_bot_5')
// (4, 8, 'sp4_r_v_b_37')
// (4, 9, 'sp4_r_v_b_24')
// (4, 10, 'sp4_r_v_b_13')
// (4, 11, 'sp4_r_v_b_0')
// (5, 6, 'neigh_op_tnl_5')
// (5, 7, 'neigh_op_lft_5')
// (5, 7, 'sp4_h_l_42')
// (5, 7, 'sp4_v_t_37')
// (5, 8, 'neigh_op_bnl_5')
// (5, 8, 'sp4_v_b_37')
// (5, 9, 'sp4_v_b_24')
// (5, 10, 'local_g0_5')
// (5, 10, 'lutff_1/in_0')
// (5, 10, 'sp4_v_b_13')
// (5, 11, 'sp4_v_b_0')

reg n52 = 0;
// (1, 8, 'sp4_r_v_b_37')
// (1, 9, 'sp4_r_v_b_24')
// (1, 10, 'sp4_r_v_b_13')
// (1, 11, 'sp4_r_v_b_0')
// (1, 12, 'sp4_r_v_b_41')
// (1, 13, 'sp4_r_v_b_28')
// (1, 14, 'neigh_op_tnr_2')
// (1, 14, 'sp4_r_v_b_17')
// (1, 15, 'neigh_op_rgt_2')
// (1, 15, 'sp4_r_v_b_4')
// (1, 16, 'neigh_op_bnr_2')
// (2, 7, 'sp4_v_t_37')
// (2, 8, 'sp4_v_b_37')
// (2, 9, 'sp4_v_b_24')
// (2, 10, 'sp4_v_b_13')
// (2, 11, 'local_g0_0')
// (2, 11, 'lutff_2/in_0')
// (2, 11, 'sp4_h_r_9')
// (2, 11, 'sp4_v_b_0')
// (2, 11, 'sp4_v_t_41')
// (2, 12, 'local_g2_1')
// (2, 12, 'lutff_1/in_0')
// (2, 12, 'sp4_v_b_41')
// (2, 13, 'local_g3_4')
// (2, 13, 'lutff_7/in_2')
// (2, 13, 'sp4_r_v_b_45')
// (2, 13, 'sp4_v_b_28')
// (2, 14, 'neigh_op_top_2')
// (2, 14, 'sp4_r_v_b_32')
// (2, 14, 'sp4_v_b_17')
// (2, 15, 'lutff_2/out')
// (2, 15, 'sp4_h_r_10')
// (2, 15, 'sp4_r_v_b_21')
// (2, 15, 'sp4_v_b_4')
// (2, 16, 'neigh_op_bot_2')
// (2, 16, 'sp4_r_v_b_8')
// (3, 11, 'sp4_h_r_20')
// (3, 12, 'sp4_h_r_8')
// (3, 12, 'sp4_v_t_45')
// (3, 13, 'sp4_v_b_45')
// (3, 14, 'neigh_op_tnl_2')
// (3, 14, 'sp4_v_b_32')
// (3, 15, 'neigh_op_lft_2')
// (3, 15, 'sp4_h_r_23')
// (3, 15, 'sp4_v_b_21')
// (3, 16, 'neigh_op_bnl_2')
// (3, 16, 'sp4_v_b_8')
// (4, 11, 'local_g2_1')
// (4, 11, 'lutff_2/in_1')
// (4, 11, 'sp4_h_r_33')
// (4, 12, 'local_g0_5')
// (4, 12, 'local_g1_5')
// (4, 12, 'lutff_1/in_0')
// (4, 12, 'lutff_2/in_0')
// (4, 12, 'lutff_3/in_0')
// (4, 12, 'sp4_h_r_21')
// (4, 15, 'local_g2_2')
// (4, 15, 'lutff_5/in_3')
// (4, 15, 'lutff_7/in_3')
// (4, 15, 'sp4_h_r_34')
// (5, 8, 'sp4_r_v_b_40')
// (5, 9, 'sp4_r_v_b_29')
// (5, 10, 'sp4_r_v_b_16')
// (5, 11, 'local_g2_4')
// (5, 11, 'local_g3_4')
// (5, 11, 'lutff_0/in_0')
// (5, 11, 'lutff_1/in_0')
// (5, 11, 'lutff_3/in_0')
// (5, 11, 'lutff_4/in_0')
// (5, 11, 'sp4_h_r_44')
// (5, 11, 'sp4_r_v_b_5')
// (5, 12, 'local_g3_4')
// (5, 12, 'local_g3_7')
// (5, 12, 'lutff_0/in_0')
// (5, 12, 'lutff_1/in_0')
// (5, 12, 'sp4_h_r_32')
// (5, 12, 'sp4_r_v_b_44')
// (5, 12, 'sp4_r_v_b_47')
// (5, 13, 'sp4_r_v_b_33')
// (5, 13, 'sp4_r_v_b_34')
// (5, 14, 'sp4_r_v_b_20')
// (5, 14, 'sp4_r_v_b_23')
// (5, 15, 'sp4_h_r_47')
// (5, 15, 'sp4_r_v_b_10')
// (5, 15, 'sp4_r_v_b_9')
// (6, 7, 'sp4_v_t_40')
// (6, 8, 'sp4_v_b_40')
// (6, 9, 'sp4_v_b_29')
// (6, 10, 'sp4_v_b_16')
// (6, 11, 'local_g0_5')
// (6, 11, 'local_g1_5')
// (6, 11, 'lutff_1/in_0')
// (6, 11, 'lutff_3/in_0')
// (6, 11, 'lutff_6/in_0')
// (6, 11, 'sp4_h_l_44')
// (6, 11, 'sp4_v_b_5')
// (6, 11, 'sp4_v_t_44')
// (6, 11, 'sp4_v_t_47')
// (6, 12, 'sp4_h_r_45')
// (6, 12, 'sp4_v_b_44')
// (6, 12, 'sp4_v_b_47')
// (6, 13, 'sp4_v_b_33')
// (6, 13, 'sp4_v_b_34')
// (6, 14, 'sp4_v_b_20')
// (6, 14, 'sp4_v_b_23')
// (6, 15, 'local_g0_2')
// (6, 15, 'lutff_4/in_2')
// (6, 15, 'sp4_h_l_47')
// (6, 15, 'sp4_v_b_10')
// (6, 15, 'sp4_v_b_9')
// (7, 12, 'sp4_h_l_45')

wire n53;
// (1, 9, 'sp12_h_r_1')
// (2, 9, 'sp12_h_r_2')
// (3, 9, 'sp12_h_r_5')
// (4, 9, 'sp12_h_r_6')
// (5, 9, 'local_g1_1')
// (5, 9, 'local_g1_4')
// (5, 9, 'lutff_0/in_2')
// (5, 9, 'lutff_2/in_3')
// (5, 9, 'lutff_4/in_3')
// (5, 9, 'sp12_h_r_9')
// (5, 9, 'sp4_h_r_4')
// (6, 9, 'sp12_h_r_10')
// (6, 9, 'sp4_h_r_17')
// (7, 8, 'neigh_op_tnr_3')
// (7, 9, 'neigh_op_rgt_3')
// (7, 9, 'sp12_h_r_13')
// (7, 9, 'sp4_h_r_28')
// (7, 10, 'neigh_op_bnr_3')
// (8, 6, 'local_g3_1')
// (8, 6, 'lutff_5/in_3')
// (8, 6, 'sp4_r_v_b_41')
// (8, 7, 'sp4_r_v_b_28')
// (8, 8, 'neigh_op_top_3')
// (8, 8, 'sp4_r_v_b_17')
// (8, 9, 'lutff_3/out')
// (8, 9, 'sp12_h_r_14')
// (8, 9, 'sp4_h_r_41')
// (8, 9, 'sp4_r_v_b_4')
// (8, 10, 'neigh_op_bot_3')
// (9, 5, 'sp4_v_t_41')
// (9, 6, 'sp4_v_b_41')
// (9, 7, 'sp4_v_b_28')
// (9, 8, 'neigh_op_tnl_3')
// (9, 8, 'sp4_v_b_17')
// (9, 9, 'neigh_op_lft_3')
// (9, 9, 'sp12_h_r_17')
// (9, 9, 'sp4_h_l_41')
// (9, 9, 'sp4_v_b_4')
// (9, 10, 'neigh_op_bnl_3')
// (10, 9, 'sp12_h_r_18')
// (11, 9, 'sp12_h_r_21')
// (12, 9, 'sp12_h_r_22')
// (13, 9, 'span12_horz_22')

reg n54 = 0;
// (1, 10, 'sp4_h_r_5')
// (2, 10, 'local_g0_0')
// (2, 10, 'lutff_6/in_0')
// (2, 10, 'sp4_h_r_16')
// (3, 7, 'neigh_op_tnr_6')
// (3, 8, 'neigh_op_rgt_6')
// (3, 9, 'neigh_op_bnr_6')
// (3, 10, 'sp4_h_r_29')
// (4, 7, 'neigh_op_top_6')
// (4, 7, 'sp4_r_v_b_40')
// (4, 8, 'lutff_6/out')
// (4, 8, 'sp4_r_v_b_29')
// (4, 9, 'neigh_op_bot_6')
// (4, 9, 'sp4_r_v_b_16')
// (4, 10, 'sp4_h_r_40')
// (4, 10, 'sp4_r_v_b_5')
// (5, 6, 'sp4_v_t_40')
// (5, 7, 'neigh_op_tnl_6')
// (5, 7, 'sp4_v_b_40')
// (5, 8, 'neigh_op_lft_6')
// (5, 8, 'sp4_v_b_29')
// (5, 9, 'neigh_op_bnl_6')
// (5, 9, 'sp4_v_b_16')
// (5, 10, 'sp4_h_l_40')
// (5, 10, 'sp4_v_b_5')

reg n55 = 0;
// (1, 11, 'neigh_op_tnr_4')
// (1, 12, 'neigh_op_rgt_4')
// (1, 13, 'neigh_op_bnr_4')
// (2, 11, 'neigh_op_top_4')
// (2, 12, 'local_g1_4')
// (2, 12, 'lutff_4/out')
// (2, 12, 'lutff_7/in_0')
// (2, 13, 'neigh_op_bot_4')
// (3, 11, 'neigh_op_tnl_4')
// (3, 12, 'neigh_op_lft_4')
// (3, 13, 'neigh_op_bnl_4')

reg n56 = 0;
// (1, 11, 'neigh_op_tnr_6')
// (1, 12, 'neigh_op_rgt_6')
// (1, 12, 'sp4_h_r_1')
// (1, 13, 'neigh_op_bnr_6')
// (2, 11, 'neigh_op_top_6')
// (2, 12, 'lutff_6/out')
// (2, 12, 'sp4_h_r_12')
// (2, 13, 'neigh_op_bot_6')
// (3, 11, 'neigh_op_tnl_6')
// (3, 12, 'neigh_op_lft_6')
// (3, 12, 'sp4_h_r_25')
// (3, 13, 'neigh_op_bnl_6')
// (4, 9, 'sp4_r_v_b_36')
// (4, 10, 'sp4_r_v_b_25')
// (4, 11, 'sp4_r_v_b_12')
// (4, 12, 'sp4_h_r_36')
// (4, 12, 'sp4_r_v_b_1')
// (5, 8, 'sp4_v_t_36')
// (5, 9, 'sp4_v_b_36')
// (5, 10, 'sp4_v_b_25')
// (5, 11, 'sp4_v_b_12')
// (5, 12, 'local_g1_1')
// (5, 12, 'lutff_5/in_3')
// (5, 12, 'sp4_h_l_36')
// (5, 12, 'sp4_v_b_1')

reg n57 = 0;
// (1, 11, 'neigh_op_tnr_7')
// (1, 12, 'neigh_op_rgt_7')
// (1, 13, 'neigh_op_bnr_7')
// (2, 11, 'neigh_op_top_7')
// (2, 12, 'local_g1_7')
// (2, 12, 'lutff_1/in_3')
// (2, 12, 'lutff_2/in_0')
// (2, 12, 'lutff_7/out')
// (2, 13, 'neigh_op_bot_7')
// (3, 11, 'neigh_op_tnl_7')
// (3, 12, 'neigh_op_lft_7')
// (3, 13, 'neigh_op_bnl_7')

reg n58 = 0;
// (1, 11, 'sp4_h_r_4')
// (1, 15, 'sp12_h_r_0')
// (2, 11, 'local_g0_1')
// (2, 11, 'lutff_2/in_1')
// (2, 11, 'sp4_h_r_17')
// (2, 12, 'local_g0_2')
// (2, 12, 'lutff_1/in_1')
// (2, 12, 'sp4_h_r_10')
// (2, 15, 'local_g1_3')
// (2, 15, 'lutff_6/in_2')
// (2, 15, 'sp12_h_r_3')
// (3, 11, 'sp4_h_r_28')
// (3, 12, 'sp4_h_r_23')
// (3, 15, 'sp12_h_r_4')
// (4, 8, 'sp4_r_v_b_41')
// (4, 9, 'sp4_r_v_b_28')
// (4, 10, 'sp4_r_v_b_17')
// (4, 10, 'sp4_r_v_b_39')
// (4, 11, 'local_g0_2')
// (4, 11, 'lutff_2/in_2')
// (4, 11, 'sp4_h_r_41')
// (4, 11, 'sp4_r_v_b_26')
// (4, 11, 'sp4_r_v_b_4')
// (4, 12, 'local_g2_2')
// (4, 12, 'local_g3_2')
// (4, 12, 'lutff_1/in_1')
// (4, 12, 'lutff_2/in_1')
// (4, 12, 'lutff_3/in_1')
// (4, 12, 'sp4_h_r_34')
// (4, 12, 'sp4_r_v_b_15')
// (4, 12, 'sp4_r_v_b_42')
// (4, 13, 'sp4_r_v_b_2')
// (4, 13, 'sp4_r_v_b_31')
// (4, 14, 'neigh_op_tnr_0')
// (4, 14, 'sp4_r_v_b_18')
// (4, 15, 'neigh_op_rgt_0')
// (4, 15, 'sp12_h_r_7')
// (4, 15, 'sp4_r_v_b_7')
// (4, 16, 'neigh_op_bnr_0')
// (5, 3, 'sp12_v_t_23')
// (5, 4, 'sp12_v_b_23')
// (5, 5, 'sp12_v_b_20')
// (5, 6, 'sp12_v_b_19')
// (5, 7, 'sp12_v_b_16')
// (5, 7, 'sp4_v_t_41')
// (5, 8, 'sp12_v_b_15')
// (5, 8, 'sp4_v_b_41')
// (5, 9, 'sp12_v_b_12')
// (5, 9, 'sp4_r_v_b_42')
// (5, 9, 'sp4_v_b_28')
// (5, 9, 'sp4_v_t_39')
// (5, 10, 'sp12_v_b_11')
// (5, 10, 'sp4_r_v_b_31')
// (5, 10, 'sp4_v_b_17')
// (5, 10, 'sp4_v_b_39')
// (5, 11, 'local_g2_0')
// (5, 11, 'local_g3_0')
// (5, 11, 'lutff_0/in_1')
// (5, 11, 'lutff_1/in_1')
// (5, 11, 'lutff_3/in_1')
// (5, 11, 'lutff_4/in_1')
// (5, 11, 'sp12_v_b_8')
// (5, 11, 'sp4_h_l_41')
// (5, 11, 'sp4_h_r_10')
// (5, 11, 'sp4_r_v_b_18')
// (5, 11, 'sp4_v_b_26')
// (5, 11, 'sp4_v_b_4')
// (5, 11, 'sp4_v_t_42')
// (5, 12, 'local_g1_7')
// (5, 12, 'local_g2_7')
// (5, 12, 'lutff_0/in_1')
// (5, 12, 'lutff_1/in_1')
// (5, 12, 'sp12_v_b_7')
// (5, 12, 'sp4_h_r_47')
// (5, 12, 'sp4_r_v_b_7')
// (5, 12, 'sp4_v_b_15')
// (5, 12, 'sp4_v_b_42')
// (5, 13, 'sp12_v_b_4')
// (5, 13, 'sp4_r_v_b_41')
// (5, 13, 'sp4_v_b_2')
// (5, 13, 'sp4_v_b_31')
// (5, 14, 'local_g0_0')
// (5, 14, 'lutff_7/in_1')
// (5, 14, 'neigh_op_top_0')
// (5, 14, 'sp12_v_b_3')
// (5, 14, 'sp4_r_v_b_28')
// (5, 14, 'sp4_v_b_18')
// (5, 15, 'lutff_0/out')
// (5, 15, 'sp12_h_r_8')
// (5, 15, 'sp12_v_b_0')
// (5, 15, 'sp4_r_v_b_17')
// (5, 15, 'sp4_v_b_7')
// (5, 16, 'neigh_op_bot_0')
// (5, 16, 'sp4_r_v_b_4')
// (6, 8, 'sp4_v_t_42')
// (6, 9, 'sp4_v_b_42')
// (6, 10, 'sp4_v_b_31')
// (6, 11, 'local_g0_2')
// (6, 11, 'local_g0_7')
// (6, 11, 'lutff_1/in_1')
// (6, 11, 'lutff_3/in_1')
// (6, 11, 'lutff_6/in_1')
// (6, 11, 'sp4_h_r_23')
// (6, 11, 'sp4_v_b_18')
// (6, 12, 'sp4_h_l_47')
// (6, 12, 'sp4_v_b_7')
// (6, 12, 'sp4_v_t_41')
// (6, 13, 'sp4_v_b_41')
// (6, 14, 'neigh_op_tnl_0')
// (6, 14, 'sp4_v_b_28')
// (6, 15, 'neigh_op_lft_0')
// (6, 15, 'sp12_h_r_11')
// (6, 15, 'sp4_v_b_17')
// (6, 16, 'neigh_op_bnl_0')
// (6, 16, 'sp4_v_b_4')
// (7, 11, 'sp4_h_r_34')
// (7, 15, 'sp12_h_r_12')
// (8, 11, 'sp4_h_r_47')
// (8, 15, 'sp12_h_r_15')
// (9, 11, 'sp4_h_l_47')
// (9, 15, 'sp12_h_r_16')
// (10, 15, 'sp12_h_r_19')
// (11, 15, 'sp12_h_r_20')
// (12, 15, 'sp12_h_r_23')
// (13, 15, 'span12_horz_23')

reg n59 = 0;
// (1, 11, 'sp4_h_r_7')
// (2, 11, 'local_g0_2')
// (2, 11, 'lutff_6/in_0')
// (2, 11, 'sp4_h_r_18')
// (3, 10, 'neigh_op_tnr_5')
// (3, 11, 'neigh_op_rgt_5')
// (3, 11, 'sp4_h_r_31')
// (3, 12, 'neigh_op_bnr_5')
// (4, 10, 'neigh_op_top_5')
// (4, 11, 'lutff_5/out')
// (4, 11, 'sp4_h_r_42')
// (4, 12, 'neigh_op_bot_5')
// (5, 10, 'neigh_op_tnl_5')
// (5, 11, 'neigh_op_lft_5')
// (5, 11, 'sp4_h_l_42')
// (5, 12, 'neigh_op_bnl_5')

reg n60 = 0;
// (1, 11, 'sp4_r_v_b_45')
// (1, 12, 'sp4_r_v_b_32')
// (1, 13, 'sp4_r_v_b_21')
// (1, 14, 'sp4_r_v_b_8')
// (2, 10, 'sp4_h_r_2')
// (2, 10, 'sp4_v_t_45')
// (2, 11, 'local_g2_5')
// (2, 11, 'lutff_2/in_3')
// (2, 11, 'sp4_v_b_45')
// (2, 12, 'sp4_v_b_32')
// (2, 13, 'sp4_v_b_21')
// (2, 14, 'sp4_v_b_8')
// (3, 9, 'neigh_op_tnr_5')
// (3, 10, 'neigh_op_rgt_5')
// (3, 10, 'sp4_h_r_15')
// (3, 11, 'neigh_op_bnr_5')
// (4, 9, 'neigh_op_top_5')
// (4, 10, 'lutff_5/out')
// (4, 10, 'sp4_h_r_26')
// (4, 11, 'neigh_op_bot_5')
// (5, 9, 'neigh_op_tnl_5')
// (5, 10, 'neigh_op_lft_5')
// (5, 10, 'sp4_h_r_39')
// (5, 11, 'neigh_op_bnl_5')
// (6, 10, 'sp4_h_l_39')

reg n61 = 0;
// (1, 12, 'sp4_r_v_b_43')
// (1, 13, 'sp4_r_v_b_30')
// (1, 14, 'sp4_r_v_b_19')
// (1, 15, 'sp4_r_v_b_6')
// (2, 11, 'sp4_h_r_0')
// (2, 11, 'sp4_v_t_43')
// (2, 12, 'local_g3_3')
// (2, 12, 'lutff_6/in_0')
// (2, 12, 'sp4_v_b_43')
// (2, 13, 'sp4_v_b_30')
// (2, 14, 'sp4_v_b_19')
// (2, 15, 'sp4_v_b_6')
// (3, 10, 'neigh_op_tnr_4')
// (3, 11, 'neigh_op_rgt_4')
// (3, 11, 'sp4_h_r_13')
// (3, 12, 'neigh_op_bnr_4')
// (4, 10, 'neigh_op_top_4')
// (4, 11, 'lutff_4/out')
// (4, 11, 'sp4_h_r_24')
// (4, 12, 'neigh_op_bot_4')
// (5, 10, 'neigh_op_tnl_4')
// (5, 11, 'neigh_op_lft_4')
// (5, 11, 'sp4_h_r_37')
// (5, 12, 'neigh_op_bnl_4')
// (6, 11, 'sp4_h_l_37')

wire n62;
// (1, 15, 'sp12_h_r_1')
// (2, 15, 'sp12_h_r_2')
// (3, 14, 'neigh_op_tnr_7')
// (3, 15, 'neigh_op_rgt_7')
// (3, 15, 'sp12_h_r_5')
// (3, 16, 'neigh_op_bnr_7')
// (4, 14, 'neigh_op_top_7')
// (4, 15, 'lutff_7/out')
// (4, 15, 'sp12_h_r_6')
// (4, 16, 'neigh_op_bot_7')
// (5, 14, 'neigh_op_tnl_7')
// (5, 15, 'local_g1_1')
// (5, 15, 'lutff_2/in_2')
// (5, 15, 'neigh_op_lft_7')
// (5, 15, 'sp12_h_r_9')
// (5, 16, 'neigh_op_bnl_7')
// (6, 15, 'sp12_h_r_10')
// (7, 15, 'sp12_h_r_13')
// (8, 15, 'sp12_h_r_14')
// (9, 15, 'sp12_h_r_17')
// (10, 15, 'sp12_h_r_18')
// (11, 15, 'sp12_h_r_21')
// (12, 15, 'sp12_h_r_22')
// (13, 15, 'span12_horz_22')

wire n63;
// (1, 15, 'sp4_h_r_5')
// (2, 15, 'local_g0_0')
// (2, 15, 'lutff_2/in_0')
// (2, 15, 'lutff_6/in_0')
// (2, 15, 'sp4_h_r_16')
// (3, 14, 'neigh_op_tnr_4')
// (3, 15, 'neigh_op_rgt_4')
// (3, 15, 'sp4_h_r_29')
// (3, 16, 'neigh_op_bnr_4')
// (4, 14, 'neigh_op_top_4')
// (4, 15, 'local_g2_4')
// (4, 15, 'lutff_0/in_2')
// (4, 15, 'lutff_4/out')
// (4, 15, 'sp4_h_r_40')
// (4, 16, 'neigh_op_bot_4')
// (5, 14, 'neigh_op_tnl_4')
// (5, 15, 'neigh_op_lft_4')
// (5, 15, 'sp4_h_l_40')
// (5, 16, 'neigh_op_bnl_4')

wire n64;
// (1, 15, 'sp4_h_r_7')
// (2, 15, 'local_g0_2')
// (2, 15, 'lutff_2/in_2')
// (2, 15, 'sp4_h_r_18')
// (3, 14, 'neigh_op_tnr_5')
// (3, 15, 'neigh_op_rgt_5')
// (3, 15, 'sp4_h_r_31')
// (3, 16, 'neigh_op_bnr_5')
// (4, 14, 'neigh_op_top_5')
// (4, 15, 'local_g2_5')
// (4, 15, 'lutff_3/in_2')
// (4, 15, 'lutff_5/out')
// (4, 15, 'sp4_h_r_42')
// (4, 16, 'neigh_op_bot_5')
// (5, 14, 'neigh_op_tnl_5')
// (5, 15, 'neigh_op_lft_5')
// (5, 15, 'sp4_h_l_42')
// (5, 16, 'neigh_op_bnl_5')

wire n65;
// (2, 3, 'sp12_h_r_0')
// (3, 3, 'sp12_h_r_3')
// (4, 3, 'sp12_h_r_4')
// (5, 2, 'neigh_op_tnr_0')
// (5, 3, 'neigh_op_rgt_0')
// (5, 3, 'sp12_h_r_7')
// (5, 4, 'neigh_op_bnr_0')
// (6, 2, 'neigh_op_top_0')
// (6, 3, 'lutff_0/out')
// (6, 3, 'sp12_h_r_8')
// (6, 4, 'neigh_op_bot_0')
// (7, 2, 'neigh_op_tnl_0')
// (7, 3, 'neigh_op_lft_0')
// (7, 3, 'sp12_h_r_11')
// (7, 4, 'neigh_op_bnl_0')
// (8, 3, 'local_g0_4')
// (8, 3, 'lutff_0/in_0')
// (8, 3, 'lutff_3/in_1')
// (8, 3, 'sp12_h_r_12')
// (9, 3, 'sp12_h_r_15')
// (10, 3, 'sp12_h_r_16')
// (11, 3, 'sp12_h_r_19')
// (12, 3, 'sp12_h_r_20')
// (13, 3, 'span12_horz_20')

reg n66 = 0;
// (2, 4, 'local_g0_2')
// (2, 4, 'lutff_0/in_0')
// (2, 4, 'sp4_h_r_10')
// (3, 3, 'neigh_op_tnr_1')
// (3, 4, 'neigh_op_rgt_1')
// (3, 4, 'sp4_h_r_23')
// (3, 5, 'neigh_op_bnr_1')
// (4, 3, 'neigh_op_top_1')
// (4, 4, 'lutff_1/out')
// (4, 4, 'sp4_h_r_34')
// (4, 5, 'neigh_op_bot_1')
// (5, 3, 'neigh_op_tnl_1')
// (5, 4, 'neigh_op_lft_1')
// (5, 4, 'sp4_h_r_47')
// (5, 5, 'neigh_op_bnl_1')
// (6, 4, 'sp4_h_l_47')

reg n67 = 0;
// (2, 4, 'sp4_r_v_b_39')
// (2, 5, 'local_g1_2')
// (2, 5, 'lutff_1/in_0')
// (2, 5, 'sp4_r_v_b_26')
// (2, 6, 'sp4_r_v_b_15')
// (2, 7, 'sp4_r_v_b_2')
// (3, 3, 'sp4_v_t_39')
// (3, 4, 'sp4_v_b_39')
// (3, 5, 'sp4_v_b_26')
// (3, 6, 'neigh_op_tnr_2')
// (3, 6, 'sp4_v_b_15')
// (3, 7, 'neigh_op_rgt_2')
// (3, 7, 'sp4_h_r_9')
// (3, 7, 'sp4_v_b_2')
// (3, 8, 'neigh_op_bnr_2')
// (4, 6, 'neigh_op_top_2')
// (4, 7, 'lutff_2/out')
// (4, 7, 'sp4_h_r_20')
// (4, 8, 'neigh_op_bot_2')
// (5, 6, 'neigh_op_tnl_2')
// (5, 7, 'neigh_op_lft_2')
// (5, 7, 'sp4_h_r_33')
// (5, 8, 'neigh_op_bnl_2')
// (6, 7, 'sp4_h_r_44')
// (7, 7, 'sp4_h_l_44')

wire n68;
// (2, 5, 'sp12_h_r_1')
// (3, 5, 'sp12_h_r_2')
// (4, 5, 'sp12_h_r_5')
// (5, 5, 'sp12_h_r_6')
// (6, 4, 'neigh_op_tnr_1')
// (6, 5, 'neigh_op_rgt_1')
// (6, 5, 'sp12_h_r_9')
// (6, 6, 'neigh_op_bnr_1')
// (7, 4, 'neigh_op_top_1')
// (7, 5, 'local_g1_2')
// (7, 5, 'lutff_0/in_3')
// (7, 5, 'lutff_1/out')
// (7, 5, 'sp12_h_r_10')
// (7, 6, 'neigh_op_bot_1')
// (8, 4, 'neigh_op_tnl_1')
// (8, 5, 'neigh_op_lft_1')
// (8, 5, 'sp12_h_r_13')
// (8, 6, 'neigh_op_bnl_1')
// (9, 5, 'sp12_h_r_14')
// (10, 5, 'sp12_h_r_17')
// (11, 5, 'sp12_h_r_18')
// (12, 5, 'sp12_h_r_21')
// (13, 5, 'span12_horz_21')

reg n69 = 0;
// (2, 6, 'sp12_h_r_1')
// (3, 6, 'sp12_h_r_2')
// (4, 6, 'sp12_h_r_5')
// (5, 6, 'sp12_h_r_6')
// (6, 6, 'sp12_h_r_9')
// (7, 6, 'sp12_h_r_10')
// (8, 5, 'neigh_op_tnr_3')
// (8, 6, 'neigh_op_rgt_3')
// (8, 6, 'sp12_h_r_13')
// (8, 7, 'neigh_op_bnr_3')
// (9, 5, 'neigh_op_top_3')
// (9, 6, 'lutff_3/out')
// (9, 6, 'sp12_h_r_14')
// (9, 7, 'neigh_op_bot_3')
// (10, 5, 'neigh_op_tnl_3')
// (10, 6, 'neigh_op_lft_3')
// (10, 6, 'sp12_h_r_17')
// (10, 7, 'neigh_op_bnl_3')
// (11, 6, 'local_g1_2')
// (11, 6, 'lutff_5/in_0')
// (11, 6, 'sp12_h_r_18')
// (12, 6, 'sp12_h_r_21')
// (13, 6, 'span12_horz_21')

reg n70 = 0;
// (2, 7, 'local_g0_0')
// (2, 7, 'lutff_0/in_2')
// (2, 7, 'sp4_h_r_0')
// (3, 7, 'sp4_h_r_13')
// (4, 7, 'neigh_op_tnr_5')
// (4, 7, 'sp4_h_r_24')
// (4, 8, 'neigh_op_rgt_5')
// (4, 9, 'neigh_op_bnr_5')
// (5, 7, 'local_g0_5')
// (5, 7, 'lutff_2/in_1')
// (5, 7, 'neigh_op_top_5')
// (5, 7, 'sp4_h_r_37')
// (5, 8, 'lutff_5/out')
// (5, 8, 'sp4_r_v_b_43')
// (5, 9, 'neigh_op_bot_5')
// (5, 9, 'sp4_r_v_b_30')
// (5, 10, 'sp4_r_v_b_19')
// (5, 11, 'sp4_r_v_b_6')
// (6, 7, 'neigh_op_tnl_5')
// (6, 7, 'sp4_h_l_37')
// (6, 7, 'sp4_v_t_43')
// (6, 8, 'neigh_op_lft_5')
// (6, 8, 'sp4_v_b_43')
// (6, 9, 'neigh_op_bnl_5')
// (6, 9, 'sp4_v_b_30')
// (6, 10, 'sp4_v_b_19')
// (6, 11, 'sp4_v_b_6')

reg n71 = 0;
// (2, 7, 'local_g0_1')
// (2, 7, 'lutff_7/in_2')
// (2, 7, 'sp4_h_r_1')
// (3, 7, 'sp4_h_r_12')
// (4, 6, 'neigh_op_tnr_2')
// (4, 7, 'neigh_op_rgt_2')
// (4, 7, 'sp4_h_r_25')
// (4, 8, 'neigh_op_bnr_2')
// (5, 6, 'neigh_op_top_2')
// (5, 7, 'local_g1_2')
// (5, 7, 'lutff_2/out')
// (5, 7, 'lutff_4/in_1')
// (5, 7, 'sp4_h_r_36')
// (5, 8, 'neigh_op_bot_2')
// (6, 6, 'neigh_op_tnl_2')
// (6, 7, 'neigh_op_lft_2')
// (6, 7, 'sp4_h_l_36')
// (6, 8, 'neigh_op_bnl_2')

reg n72 = 0;
// (2, 7, 'sp12_h_r_0')
// (3, 7, 'sp12_h_r_3')
// (4, 7, 'sp12_h_r_4')
// (5, 7, 'sp12_h_r_7')
// (6, 7, 'sp12_h_r_8')
// (7, 6, 'neigh_op_tnr_2')
// (7, 7, 'neigh_op_rgt_2')
// (7, 7, 'sp12_h_r_11')
// (7, 8, 'neigh_op_bnr_2')
// (8, 6, 'neigh_op_top_2')
// (8, 7, 'local_g0_2')
// (8, 7, 'lutff_2/out')
// (8, 7, 'lutff_7/in_1')
// (8, 7, 'sp12_h_r_12')
// (8, 8, 'neigh_op_bot_2')
// (9, 6, 'neigh_op_tnl_2')
// (9, 7, 'neigh_op_lft_2')
// (9, 7, 'sp12_h_r_15')
// (9, 8, 'neigh_op_bnl_2')
// (10, 7, 'sp12_h_r_16')
// (11, 7, 'local_g1_3')
// (11, 7, 'lutff_0/in_2')
// (11, 7, 'sp12_h_r_19')
// (12, 7, 'sp12_h_r_20')
// (13, 7, 'span12_horz_20')

reg n73 = 0;
// (2, 7, 'sp12_h_r_1')
// (3, 7, 'sp12_h_r_2')
// (4, 7, 'sp12_h_r_5')
// (5, 7, 'sp12_h_r_6')
// (6, 7, 'sp12_h_r_9')
// (7, 7, 'sp12_h_r_10')
// (8, 6, 'neigh_op_tnr_3')
// (8, 7, 'neigh_op_rgt_3')
// (8, 7, 'sp12_h_r_13')
// (8, 8, 'neigh_op_bnr_3')
// (9, 6, 'neigh_op_top_3')
// (9, 7, 'lutff_3/out')
// (9, 7, 'sp12_h_r_14')
// (9, 8, 'neigh_op_bot_3')
// (10, 6, 'neigh_op_tnl_3')
// (10, 7, 'neigh_op_lft_3')
// (10, 7, 'sp12_h_r_17')
// (10, 8, 'neigh_op_bnl_3')
// (11, 7, 'sp12_h_r_18')
// (12, 7, 'local_g0_5')
// (12, 7, 'lutff_1/in_0')
// (12, 7, 'sp12_h_r_21')
// (13, 7, 'span12_horz_21')

wire n74;
// (2, 12, 'sp4_h_r_0')
// (3, 11, 'neigh_op_tnr_4')
// (3, 12, 'neigh_op_rgt_4')
// (3, 12, 'sp4_h_r_13')
// (3, 13, 'neigh_op_bnr_4')
// (4, 11, 'neigh_op_top_4')
// (4, 12, 'lutff_4/out')
// (4, 12, 'sp4_h_r_24')
// (4, 13, 'neigh_op_bot_4')
// (5, 11, 'neigh_op_tnl_4')
// (5, 12, 'neigh_op_lft_4')
// (5, 12, 'sp4_h_r_37')
// (5, 13, 'neigh_op_bnl_4')
// (5, 13, 'sp4_r_v_b_37')
// (5, 14, 'sp4_r_v_b_24')
// (5, 15, 'sp4_r_v_b_13')
// (5, 16, 'sp4_r_v_b_0')
// (6, 12, 'sp4_h_l_37')
// (6, 12, 'sp4_v_t_37')
// (6, 13, 'local_g2_5')
// (6, 13, 'local_g3_5')
// (6, 13, 'lutff_2/in_3')
// (6, 13, 'lutff_3/in_1')
// (6, 13, 'lutff_5/in_2')
// (6, 13, 'lutff_7/in_2')
// (6, 13, 'sp4_v_b_37')
// (6, 14, 'sp4_v_b_24')
// (6, 15, 'sp4_v_b_13')
// (6, 16, 'sp4_v_b_0')

wire n75;
// (2, 12, 'sp4_h_r_2')
// (3, 11, 'neigh_op_tnr_5')
// (3, 12, 'neigh_op_rgt_5')
// (3, 12, 'sp4_h_r_15')
// (3, 13, 'neigh_op_bnr_5')
// (4, 11, 'neigh_op_top_5')
// (4, 12, 'lutff_5/out')
// (4, 12, 'sp4_h_r_10')
// (4, 12, 'sp4_h_r_26')
// (4, 13, 'neigh_op_bot_5')
// (5, 11, 'neigh_op_tnl_5')
// (5, 12, 'neigh_op_lft_5')
// (5, 12, 'sp4_h_r_23')
// (5, 12, 'sp4_h_r_39')
// (5, 13, 'neigh_op_bnl_5')
// (5, 13, 'sp4_r_v_b_39')
// (5, 14, 'sp4_r_v_b_26')
// (5, 15, 'sp4_r_v_b_15')
// (5, 16, 'sp4_r_v_b_2')
// (6, 12, 'local_g2_2')
// (6, 12, 'lutff_6/in_2')
// (6, 12, 'sp4_h_l_39')
// (6, 12, 'sp4_h_r_34')
// (6, 12, 'sp4_v_t_39')
// (6, 13, 'local_g2_7')
// (6, 13, 'lutff_0/in_3')
// (6, 13, 'lutff_3/in_2')
// (6, 13, 'sp4_v_b_39')
// (6, 14, 'sp4_v_b_26')
// (6, 15, 'sp4_v_b_15')
// (6, 16, 'sp4_v_b_2')
// (7, 12, 'sp4_h_r_47')
// (8, 12, 'sp4_h_l_47')

reg n76 = 0;
// (2, 13, 'sp12_h_r_1')
// (3, 13, 'sp12_h_r_2')
// (4, 13, 'sp12_h_r_5')
// (5, 13, 'sp12_h_r_6')
// (6, 13, 'sp12_h_r_9')
// (7, 13, 'sp12_h_r_10')
// (8, 12, 'neigh_op_tnr_3')
// (8, 13, 'neigh_op_rgt_3')
// (8, 13, 'sp12_h_r_13')
// (8, 13, 'sp4_h_r_6')
// (8, 14, 'neigh_op_bnr_3')
// (9, 12, 'neigh_op_top_3')
// (9, 13, 'local_g1_3')
// (9, 13, 'lutff_3/in_3')
// (9, 13, 'lutff_3/out')
// (9, 13, 'lutff_5/in_3')
// (9, 13, 'sp12_h_r_14')
// (9, 13, 'sp4_h_r_19')
// (9, 14, 'neigh_op_bot_3')
// (10, 12, 'neigh_op_tnl_3')
// (10, 13, 'neigh_op_lft_3')
// (10, 13, 'sp12_h_r_17')
// (10, 13, 'sp4_h_r_30')
// (10, 14, 'neigh_op_bnl_3')
// (11, 10, 'sp4_r_v_b_43')
// (11, 11, 'local_g0_6')
// (11, 11, 'local_g1_6')
// (11, 11, 'lutff_0/in_3')
// (11, 11, 'lutff_4/in_3')
// (11, 11, 'lutff_7/in_3')
// (11, 11, 'sp4_r_v_b_30')
// (11, 12, 'local_g3_3')
// (11, 12, 'lutff_4/in_2')
// (11, 12, 'sp4_r_v_b_19')
// (11, 13, 'local_g1_2')
// (11, 13, 'lutff_0/in_1')
// (11, 13, 'sp12_h_r_18')
// (11, 13, 'sp4_h_r_43')
// (11, 13, 'sp4_r_v_b_6')
// (12, 9, 'sp4_v_t_43')
// (12, 10, 'sp4_v_b_43')
// (12, 11, 'sp4_v_b_30')
// (12, 12, 'sp4_v_b_19')
// (12, 13, 'sp12_h_r_21')
// (12, 13, 'sp4_h_l_43')
// (12, 13, 'sp4_v_b_6')
// (13, 13, 'span12_horz_21')

wire n77;
// (2, 14, 'sp4_h_r_0')
// (3, 14, 'sp4_h_r_13')
// (4, 14, 'sp4_h_r_24')
// (5, 11, 'neigh_op_tnr_4')
// (5, 11, 'sp4_r_v_b_37')
// (5, 12, 'neigh_op_rgt_4')
// (5, 12, 'sp4_r_v_b_24')
// (5, 13, 'neigh_op_bnr_4')
// (5, 13, 'sp4_r_v_b_13')
// (5, 14, 'sp4_h_r_37')
// (5, 14, 'sp4_r_v_b_0')
// (6, 10, 'sp4_v_t_37')
// (6, 11, 'neigh_op_top_4')
// (6, 11, 'sp4_v_b_37')
// (6, 12, 'lutff_4/out')
// (6, 12, 'sp4_v_b_24')
// (6, 13, 'neigh_op_bot_4')
// (6, 13, 'sp4_v_b_13')
// (6, 14, 'local_g0_0')
// (6, 14, 'lutff_0/in_0')
// (6, 14, 'lutff_6/in_2')
// (6, 14, 'sp4_h_l_37')
// (6, 14, 'sp4_h_r_3')
// (6, 14, 'sp4_v_b_0')
// (7, 11, 'neigh_op_tnl_4')
// (7, 12, 'neigh_op_lft_4')
// (7, 13, 'neigh_op_bnl_4')
// (7, 14, 'sp4_h_r_14')
// (8, 14, 'local_g2_3')
// (8, 14, 'local_g3_3')
// (8, 14, 'lutff_3/in_3')
// (8, 14, 'lutff_4/in_2')
// (8, 14, 'lutff_7/in_2')
// (8, 14, 'sp4_h_r_27')
// (9, 14, 'sp4_h_r_38')
// (10, 14, 'sp4_h_l_38')

reg \d_out[6] = 0 ;
// (3, 1, 'sp4_r_v_b_26')
// (3, 2, 'neigh_op_tnr_1')
// (3, 2, 'sp4_r_v_b_15')
// (3, 3, 'neigh_op_rgt_1')
// (3, 3, 'sp4_r_v_b_2')
// (3, 4, 'neigh_op_bnr_1')
// (4, 0, 'io_1/D_OUT_0')
// (4, 0, 'io_1/PAD')
// (4, 0, 'local_g1_2')
// (4, 0, 'span4_vert_26')
// (4, 1, 'sp4_v_b_26')
// (4, 2, 'neigh_op_top_1')
// (4, 2, 'sp4_v_b_15')
// (4, 3, 'lutff_1/out')
// (4, 3, 'sp4_v_b_2')
// (4, 4, 'neigh_op_bot_1')
// (5, 2, 'neigh_op_tnl_1')
// (5, 3, 'neigh_op_lft_1')
// (5, 4, 'neigh_op_bnl_1')

reg n79 = 0;
// (3, 2, 'neigh_op_tnr_0')
// (3, 3, 'neigh_op_rgt_0')
// (3, 4, 'neigh_op_bnr_0')
// (4, 2, 'neigh_op_top_0')
// (4, 3, 'local_g1_0')
// (4, 3, 'lutff_0/out')
// (4, 3, 'lutff_7/in_0')
// (4, 4, 'neigh_op_bot_0')
// (5, 2, 'neigh_op_tnl_0')
// (5, 3, 'neigh_op_lft_0')
// (5, 4, 'neigh_op_bnl_0')

reg n80 = 0;
// (3, 2, 'neigh_op_tnr_3')
// (3, 3, 'neigh_op_rgt_3')
// (3, 4, 'neigh_op_bnr_3')
// (4, 2, 'neigh_op_top_3')
// (4, 3, 'local_g1_3')
// (4, 3, 'lutff_2/in_0')
// (4, 3, 'lutff_3/out')
// (4, 4, 'neigh_op_bot_3')
// (5, 2, 'neigh_op_tnl_3')
// (5, 3, 'neigh_op_lft_3')
// (5, 4, 'neigh_op_bnl_3')

reg n81 = 0;
// (3, 2, 'neigh_op_tnr_4')
// (3, 3, 'neigh_op_rgt_4')
// (3, 4, 'neigh_op_bnr_4')
// (4, 2, 'neigh_op_top_4')
// (4, 3, 'local_g0_4')
// (4, 3, 'lutff_0/in_0')
// (4, 3, 'lutff_4/out')
// (4, 4, 'neigh_op_bot_4')
// (5, 2, 'neigh_op_tnl_4')
// (5, 3, 'neigh_op_lft_4')
// (5, 4, 'neigh_op_bnl_4')

reg n82 = 0;
// (3, 2, 'neigh_op_tnr_7')
// (3, 3, 'neigh_op_rgt_7')
// (3, 4, 'neigh_op_bnr_7')
// (4, 2, 'neigh_op_top_7')
// (4, 3, 'local_g0_7')
// (4, 3, 'lutff_3/in_0')
// (4, 3, 'lutff_7/out')
// (4, 4, 'neigh_op_bot_7')
// (5, 2, 'neigh_op_tnl_7')
// (5, 3, 'neigh_op_lft_7')
// (5, 4, 'neigh_op_bnl_7')

wire n83;
// (3, 2, 'sp4_r_v_b_41')
// (3, 3, 'sp4_r_v_b_28')
// (3, 4, 'sp4_r_v_b_17')
// (3, 5, 'sp4_r_v_b_4')
// (3, 6, 'sp4_r_v_b_36')
// (3, 7, 'sp4_r_v_b_25')
// (3, 8, 'sp4_r_v_b_12')
// (3, 9, 'sp4_r_v_b_1')
// (4, 1, 'sp4_v_t_41')
// (4, 2, 'sp4_r_v_b_41')
// (4, 2, 'sp4_v_b_41')
// (4, 3, 'sp4_r_v_b_28')
// (4, 3, 'sp4_v_b_28')
// (4, 4, 'local_g0_1')
// (4, 4, 'lutff_1/in_2')
// (4, 4, 'sp4_r_v_b_17')
// (4, 4, 'sp4_v_b_17')
// (4, 5, 'sp4_r_v_b_4')
// (4, 5, 'sp4_v_b_4')
// (4, 5, 'sp4_v_t_36')
// (4, 6, 'sp4_r_v_b_36')
// (4, 6, 'sp4_v_b_36')
// (4, 7, 'sp4_r_v_b_25')
// (4, 7, 'sp4_v_b_25')
// (4, 8, 'sp4_r_v_b_12')
// (4, 8, 'sp4_v_b_12')
// (4, 9, 'sp4_h_r_8')
// (4, 9, 'sp4_r_v_b_1')
// (4, 9, 'sp4_v_b_1')
// (4, 10, 'sp4_r_v_b_40')
// (4, 11, 'sp4_r_v_b_29')
// (4, 12, 'sp4_r_v_b_16')
// (4, 13, 'sp4_r_v_b_5')
// (5, 1, 'sp4_v_t_41')
// (5, 2, 'sp4_v_b_41')
// (5, 3, 'sp4_v_b_28')
// (5, 4, 'local_g0_1')
// (5, 4, 'lutff_0/in_1')
// (5, 4, 'lutff_4/in_1')
// (5, 4, 'sp4_v_b_17')
// (5, 5, 'sp4_v_b_4')
// (5, 5, 'sp4_v_t_36')
// (5, 6, 'sp4_v_b_36')
// (5, 7, 'sp4_v_b_25')
// (5, 8, 'sp4_v_b_12')
// (5, 9, 'sp4_h_r_21')
// (5, 9, 'sp4_v_b_1')
// (5, 9, 'sp4_v_t_40')
// (5, 10, 'sp4_v_b_40')
// (5, 11, 'sp4_v_b_29')
// (5, 12, 'sp4_v_b_16')
// (5, 13, 'sp4_h_r_5')
// (5, 13, 'sp4_v_b_5')
// (6, 9, 'sp4_h_r_32')
// (6, 13, 'sp4_h_r_16')
// (7, 9, 'sp4_h_r_45')
// (7, 10, 'sp4_r_v_b_45')
// (7, 11, 'sp4_r_v_b_32')
// (7, 12, 'neigh_op_tnr_4')
// (7, 12, 'sp4_r_v_b_21')
// (7, 13, 'neigh_op_rgt_4')
// (7, 13, 'sp4_h_r_29')
// (7, 13, 'sp4_r_v_b_8')
// (7, 14, 'neigh_op_bnr_4')
// (8, 9, 'sp4_h_l_45')
// (8, 9, 'sp4_v_t_45')
// (8, 10, 'sp4_v_b_45')
// (8, 11, 'sp4_v_b_32')
// (8, 12, 'neigh_op_top_4')
// (8, 12, 'sp4_v_b_21')
// (8, 13, 'lutff_4/out')
// (8, 13, 'sp4_h_r_40')
// (8, 13, 'sp4_v_b_8')
// (8, 14, 'neigh_op_bot_4')
// (9, 12, 'neigh_op_tnl_4')
// (9, 13, 'neigh_op_lft_4')
// (9, 13, 'sp4_h_l_40')
// (9, 14, 'neigh_op_bnl_4')

wire n84;
// (3, 4, 'sp4_h_r_9')
// (3, 6, 'sp4_h_r_4')
// (4, 4, 'sp4_h_r_20')
// (4, 6, 'local_g0_1')
// (4, 6, 'lutff_1/in_2')
// (4, 6, 'sp4_h_r_17')
// (5, 4, 'local_g2_1')
// (5, 4, 'lutff_2/in_1')
// (5, 4, 'sp4_h_r_33')
// (5, 6, 'sp4_h_r_28')
// (6, 3, 'sp4_r_v_b_46')
// (6, 4, 'local_g0_0')
// (6, 4, 'lutff_7/in_1')
// (6, 4, 'sp4_h_r_44')
// (6, 4, 'sp4_r_v_b_35')
// (6, 5, 'sp4_r_v_b_22')
// (6, 5, 'sp4_r_v_b_44')
// (6, 6, 'sp4_h_r_41')
// (6, 6, 'sp4_r_v_b_11')
// (6, 6, 'sp4_r_v_b_33')
// (6, 7, 'sp4_r_v_b_20')
// (6, 8, 'sp4_r_v_b_9')
// (6, 11, 'neigh_op_tnr_3')
// (6, 12, 'neigh_op_rgt_3')
// (6, 13, 'neigh_op_bnr_3')
// (7, 2, 'sp4_v_t_46')
// (7, 3, 'sp12_v_t_22')
// (7, 3, 'sp4_v_b_46')
// (7, 4, 'sp12_v_b_22')
// (7, 4, 'sp4_h_l_44')
// (7, 4, 'sp4_v_b_35')
// (7, 4, 'sp4_v_t_44')
// (7, 5, 'sp12_v_b_21')
// (7, 5, 'sp4_v_b_22')
// (7, 5, 'sp4_v_b_44')
// (7, 6, 'sp12_v_b_18')
// (7, 6, 'sp4_h_l_41')
// (7, 6, 'sp4_v_b_11')
// (7, 6, 'sp4_v_b_33')
// (7, 7, 'sp12_v_b_17')
// (7, 7, 'sp4_v_b_20')
// (7, 8, 'sp12_v_b_14')
// (7, 8, 'sp4_v_b_9')
// (7, 9, 'sp12_v_b_13')
// (7, 10, 'sp12_v_b_10')
// (7, 11, 'neigh_op_top_3')
// (7, 11, 'sp12_v_b_9')
// (7, 12, 'lutff_3/out')
// (7, 12, 'sp12_v_b_6')
// (7, 13, 'neigh_op_bot_3')
// (7, 13, 'sp12_v_b_5')
// (7, 14, 'sp12_v_b_2')
// (7, 15, 'sp12_v_b_1')
// (8, 11, 'neigh_op_tnl_3')
// (8, 12, 'neigh_op_lft_3')
// (8, 13, 'neigh_op_bnl_3')

reg n85 = 0;
// (3, 4, 'sp4_r_v_b_38')
// (3, 5, 'neigh_op_tnr_7')
// (3, 5, 'sp4_r_v_b_27')
// (3, 6, 'neigh_op_rgt_7')
// (3, 6, 'sp4_r_v_b_14')
// (3, 7, 'neigh_op_bnr_7')
// (3, 7, 'sp4_r_v_b_3')
// (4, 3, 'sp4_v_t_38')
// (4, 4, 'sp4_v_b_38')
// (4, 5, 'neigh_op_top_7')
// (4, 5, 'sp4_v_b_27')
// (4, 6, 'lutff_7/out')
// (4, 6, 'sp4_v_b_14')
// (4, 7, 'local_g0_3')
// (4, 7, 'lutff_5/in_0')
// (4, 7, 'neigh_op_bot_7')
// (4, 7, 'sp4_v_b_3')
// (5, 5, 'neigh_op_tnl_7')
// (5, 6, 'neigh_op_lft_7')
// (5, 7, 'neigh_op_bnl_7')

reg n86 = 0;
// (3, 5, 'neigh_op_tnr_1')
// (3, 6, 'neigh_op_rgt_1')
// (3, 7, 'neigh_op_bnr_1')
// (4, 5, 'neigh_op_top_1')
// (4, 6, 'lutff_1/out')
// (4, 7, 'local_g0_1')
// (4, 7, 'lutff_7/in_0')
// (4, 7, 'neigh_op_bot_1')
// (5, 5, 'neigh_op_tnl_1')
// (5, 6, 'neigh_op_lft_1')
// (5, 7, 'neigh_op_bnl_1')

reg n87 = 0;
// (3, 5, 'neigh_op_tnr_3')
// (3, 6, 'neigh_op_rgt_3')
// (3, 7, 'neigh_op_bnr_3')
// (4, 5, 'neigh_op_top_3')
// (4, 6, 'lutff_3/out')
// (4, 7, 'local_g1_3')
// (4, 7, 'lutff_0/in_0')
// (4, 7, 'neigh_op_bot_3')
// (5, 5, 'neigh_op_tnl_3')
// (5, 6, 'neigh_op_lft_3')
// (5, 7, 'neigh_op_bnl_3')

wire n88;
// (3, 5, 'sp4_r_v_b_36')
// (3, 6, 'sp4_r_v_b_25')
// (3, 7, 'sp4_r_v_b_12')
// (3, 8, 'sp4_r_v_b_1')
// (4, 4, 'sp4_v_t_36')
// (4, 5, 'sp4_v_b_36')
// (4, 6, 'local_g2_1')
// (4, 6, 'lutff_3/in_0')
// (4, 6, 'sp4_v_b_25')
// (4, 7, 'sp4_v_b_12')
// (4, 8, 'sp4_h_r_8')
// (4, 8, 'sp4_v_b_1')
// (5, 8, 'sp4_h_r_21')
// (6, 8, 'sp4_h_r_32')
// (7, 5, 'sp4_r_v_b_38')
// (7, 6, 'sp4_r_v_b_27')
// (7, 7, 'sp4_r_v_b_14')
// (7, 8, 'sp4_h_r_45')
// (7, 8, 'sp4_r_v_b_3')
// (7, 9, 'sp4_r_v_b_37')
// (7, 10, 'sp4_r_v_b_24')
// (7, 11, 'neigh_op_tnr_0')
// (7, 11, 'sp4_r_v_b_13')
// (7, 12, 'neigh_op_rgt_0')
// (7, 12, 'sp4_r_v_b_0')
// (7, 13, 'neigh_op_bnr_0')
// (8, 4, 'sp4_v_t_38')
// (8, 5, 'sp4_v_b_38')
// (8, 6, 'local_g2_3')
// (8, 6, 'local_g3_3')
// (8, 6, 'lutff_5/in_2')
// (8, 6, 'lutff_6/in_2')
// (8, 6, 'sp4_v_b_27')
// (8, 7, 'sp4_v_b_14')
// (8, 8, 'sp4_h_l_45')
// (8, 8, 'sp4_v_b_3')
// (8, 8, 'sp4_v_t_37')
// (8, 9, 'sp4_v_b_37')
// (8, 10, 'sp4_v_b_24')
// (8, 11, 'neigh_op_top_0')
// (8, 11, 'sp4_v_b_13')
// (8, 12, 'lutff_0/out')
// (8, 12, 'sp4_v_b_0')
// (8, 13, 'neigh_op_bot_0')
// (9, 11, 'neigh_op_tnl_0')
// (9, 12, 'neigh_op_lft_0')
// (9, 13, 'neigh_op_bnl_0')

reg n89 = 0;
// (3, 6, 'neigh_op_tnr_0')
// (3, 7, 'neigh_op_rgt_0')
// (3, 8, 'neigh_op_bnr_0')
// (4, 6, 'neigh_op_top_0')
// (4, 7, 'lutff_0/out')
// (4, 8, 'neigh_op_bot_0')
// (5, 6, 'neigh_op_tnl_0')
// (5, 7, 'local_g1_0')
// (5, 7, 'lutff_5/in_0')
// (5, 7, 'neigh_op_lft_0')
// (5, 8, 'neigh_op_bnl_0')

reg n90 = 0;
// (3, 6, 'neigh_op_tnr_1')
// (3, 7, 'neigh_op_rgt_1')
// (3, 7, 'sp4_h_r_7')
// (3, 8, 'neigh_op_bnr_1')
// (4, 4, 'sp12_v_t_22')
// (4, 4, 'sp4_r_v_b_38')
// (4, 5, 'sp12_v_b_22')
// (4, 5, 'sp4_r_v_b_27')
// (4, 6, 'neigh_op_top_1')
// (4, 6, 'sp12_v_b_21')
// (4, 6, 'sp4_r_v_b_14')
// (4, 7, 'lutff_1/out')
// (4, 7, 'sp12_v_b_18')
// (4, 7, 'sp4_h_r_18')
// (4, 7, 'sp4_r_v_b_3')
// (4, 8, 'neigh_op_bot_1')
// (4, 8, 'sp12_v_b_17')
// (4, 9, 'sp12_v_b_14')
// (4, 10, 'sp12_v_b_13')
// (4, 11, 'sp12_v_b_10')
// (4, 12, 'local_g3_1')
// (4, 12, 'lutff_6/in_0')
// (4, 12, 'sp12_v_b_9')
// (4, 13, 'sp12_v_b_6')
// (4, 14, 'sp12_v_b_5')
// (4, 15, 'sp12_v_b_2')
// (4, 16, 'sp12_v_b_1')
// (5, 3, 'sp4_v_t_38')
// (5, 4, 'sp4_v_b_38')
// (5, 5, 'local_g3_3')
// (5, 5, 'lutff_2/in_0')
// (5, 5, 'sp4_v_b_27')
// (5, 6, 'neigh_op_tnl_1')
// (5, 6, 'sp4_v_b_14')
// (5, 7, 'neigh_op_lft_1')
// (5, 7, 'sp4_h_r_31')
// (5, 7, 'sp4_v_b_3')
// (5, 8, 'neigh_op_bnl_1')
// (6, 4, 'sp4_r_v_b_36')
// (6, 5, 'sp4_r_v_b_25')
// (6, 6, 'local_g2_4')
// (6, 6, 'lutff_1/in_3')
// (6, 6, 'sp4_r_v_b_12')
// (6, 7, 'sp4_h_r_42')
// (6, 7, 'sp4_r_v_b_1')
// (7, 3, 'sp4_v_t_36')
// (7, 4, 'sp4_v_b_36')
// (7, 5, 'sp4_v_b_25')
// (7, 6, 'sp4_v_b_12')
// (7, 7, 'sp4_h_l_42')
// (7, 7, 'sp4_v_b_1')

reg n91 = 0;
// (3, 6, 'neigh_op_tnr_3')
// (3, 7, 'neigh_op_rgt_3')
// (3, 7, 'sp4_r_v_b_38')
// (3, 8, 'neigh_op_bnr_3')
// (3, 8, 'sp4_r_v_b_27')
// (3, 9, 'sp4_r_v_b_14')
// (3, 10, 'sp4_r_v_b_3')
// (4, 5, 'sp4_r_v_b_47')
// (4, 6, 'neigh_op_top_3')
// (4, 6, 'sp4_r_v_b_34')
// (4, 6, 'sp4_v_t_38')
// (4, 7, 'lutff_3/out')
// (4, 7, 'sp4_r_v_b_23')
// (4, 7, 'sp4_v_b_38')
// (4, 8, 'neigh_op_bot_3')
// (4, 8, 'sp4_r_v_b_10')
// (4, 8, 'sp4_v_b_27')
// (4, 9, 'sp4_r_v_b_47')
// (4, 9, 'sp4_v_b_14')
// (4, 10, 'sp4_h_r_9')
// (4, 10, 'sp4_r_v_b_34')
// (4, 10, 'sp4_v_b_3')
// (4, 11, 'sp4_r_v_b_23')
// (4, 12, 'sp4_r_v_b_10')
// (5, 4, 'sp4_v_t_47')
// (5, 5, 'sp4_v_b_47')
// (5, 6, 'neigh_op_tnl_3')
// (5, 6, 'sp4_v_b_34')
// (5, 7, 'neigh_op_lft_3')
// (5, 7, 'sp4_v_b_23')
// (5, 8, 'neigh_op_bnl_3')
// (5, 8, 'sp4_v_b_10')
// (5, 8, 'sp4_v_t_47')
// (5, 9, 'sp4_v_b_47')
// (5, 10, 'local_g0_4')
// (5, 10, 'lutff_2/in_0')
// (5, 10, 'sp4_h_r_20')
// (5, 10, 'sp4_v_b_34')
// (5, 11, 'sp4_v_b_23')
// (5, 12, 'local_g0_2')
// (5, 12, 'lutff_1/in_3')
// (5, 12, 'sp4_v_b_10')
// (6, 10, 'sp4_h_r_33')
// (7, 10, 'sp4_h_r_44')
// (8, 10, 'sp4_h_l_44')

reg n92 = 0;
// (3, 6, 'neigh_op_tnr_6')
// (3, 7, 'neigh_op_rgt_6')
// (3, 8, 'neigh_op_bnr_6')
// (4, 6, 'neigh_op_top_6')
// (4, 7, 'local_g0_6')
// (4, 7, 'lutff_2/in_0')
// (4, 7, 'lutff_6/out')
// (4, 8, 'neigh_op_bot_6')
// (5, 6, 'neigh_op_tnl_6')
// (5, 7, 'neigh_op_lft_6')
// (5, 8, 'neigh_op_bnl_6')

reg n93 = 0;
// (3, 6, 'neigh_op_tnr_7')
// (3, 7, 'neigh_op_rgt_7')
// (3, 8, 'neigh_op_bnr_7')
// (4, 6, 'neigh_op_top_7')
// (4, 7, 'local_g0_7')
// (4, 7, 'lutff_3/in_0')
// (4, 7, 'lutff_7/out')
// (4, 8, 'neigh_op_bot_7')
// (5, 6, 'neigh_op_tnl_7')
// (5, 7, 'neigh_op_lft_7')
// (5, 8, 'neigh_op_bnl_7')

reg n94 = 0;
// (3, 7, 'neigh_op_tnr_0')
// (3, 8, 'neigh_op_rgt_0')
// (3, 9, 'neigh_op_bnr_0')
// (4, 7, 'neigh_op_top_0')
// (4, 8, 'local_g1_0')
// (4, 8, 'lutff_0/out')
// (4, 8, 'lutff_1/in_0')
// (4, 9, 'neigh_op_bot_0')
// (5, 7, 'neigh_op_tnl_0')
// (5, 8, 'neigh_op_lft_0')
// (5, 9, 'neigh_op_bnl_0')

reg n95 = 0;
// (3, 7, 'neigh_op_tnr_1')
// (3, 8, 'neigh_op_rgt_1')
// (3, 9, 'neigh_op_bnr_1')
// (4, 7, 'neigh_op_top_1')
// (4, 8, 'local_g1_1')
// (4, 8, 'lutff_1/out')
// (4, 8, 'lutff_6/in_0')
// (4, 9, 'neigh_op_bot_1')
// (5, 7, 'neigh_op_tnl_1')
// (5, 8, 'neigh_op_lft_1')
// (5, 9, 'neigh_op_bnl_1')

reg n96 = 0;
// (3, 7, 'neigh_op_tnr_2')
// (3, 8, 'neigh_op_rgt_2')
// (3, 9, 'neigh_op_bnr_2')
// (4, 7, 'neigh_op_top_2')
// (4, 8, 'lutff_2/out')
// (4, 9, 'neigh_op_bot_2')
// (5, 7, 'neigh_op_tnl_2')
// (5, 8, 'local_g0_2')
// (5, 8, 'lutff_0/in_0')
// (5, 8, 'neigh_op_lft_2')
// (5, 9, 'neigh_op_bnl_2')

reg n97 = 0;
// (3, 7, 'neigh_op_tnr_3')
// (3, 8, 'neigh_op_rgt_3')
// (3, 9, 'neigh_op_bnr_3')
// (4, 7, 'neigh_op_top_3')
// (4, 8, 'local_g1_3')
// (4, 8, 'lutff_0/in_0')
// (4, 8, 'lutff_3/out')
// (4, 9, 'neigh_op_bot_3')
// (5, 7, 'neigh_op_tnl_3')
// (5, 8, 'neigh_op_lft_3')
// (5, 9, 'neigh_op_bnl_3')

reg \d_out[7] = 0 ;
// (3, 7, 'neigh_op_tnr_4')
// (3, 8, 'neigh_op_rgt_4')
// (3, 9, 'neigh_op_bnr_4')
// (4, 0, 'io_0/D_OUT_0')
// (4, 0, 'io_0/PAD')
// (4, 0, 'local_g1_7')
// (4, 0, 'span12_vert_23')
// (4, 1, 'sp12_v_b_23')
// (4, 2, 'sp12_v_b_20')
// (4, 3, 'sp12_v_b_19')
// (4, 4, 'sp12_v_b_16')
// (4, 5, 'sp12_v_b_15')
// (4, 6, 'sp12_v_b_12')
// (4, 7, 'neigh_op_top_4')
// (4, 7, 'sp12_v_b_11')
// (4, 8, 'lutff_4/out')
// (4, 8, 'sp12_v_b_8')
// (4, 9, 'neigh_op_bot_4')
// (4, 9, 'sp12_v_b_7')
// (4, 10, 'sp12_v_b_4')
// (4, 11, 'sp12_v_b_3')
// (4, 12, 'sp12_v_b_0')
// (5, 7, 'neigh_op_tnl_4')
// (5, 8, 'neigh_op_lft_4')
// (5, 9, 'neigh_op_bnl_4')

reg n99 = 0;
// (3, 7, 'neigh_op_tnr_5')
// (3, 8, 'neigh_op_rgt_5')
// (3, 9, 'neigh_op_bnr_5')
// (4, 7, 'neigh_op_top_5')
// (4, 8, 'local_g2_5')
// (4, 8, 'lutff_3/in_0')
// (4, 8, 'lutff_5/out')
// (4, 9, 'neigh_op_bot_5')
// (5, 7, 'neigh_op_tnl_5')
// (5, 8, 'neigh_op_lft_5')
// (5, 9, 'neigh_op_bnl_5')

reg n100 = 0;
// (3, 7, 'neigh_op_tnr_7')
// (3, 8, 'neigh_op_rgt_7')
// (3, 9, 'neigh_op_bnr_7')
// (4, 7, 'neigh_op_top_7')
// (4, 8, 'local_g1_7')
// (4, 8, 'lutff_2/in_0')
// (4, 8, 'lutff_7/out')
// (4, 9, 'neigh_op_bot_7')
// (5, 7, 'neigh_op_tnl_7')
// (5, 8, 'neigh_op_lft_7')
// (5, 9, 'neigh_op_bnl_7')

wire n101;
// (3, 7, 'sp4_h_r_11')
// (4, 7, 'sp4_h_r_22')
// (5, 7, 'sp4_h_r_35')
// (6, 4, 'sp4_r_v_b_40')
// (6, 5, 'sp4_r_v_b_29')
// (6, 6, 'sp4_r_v_b_16')
// (6, 7, 'local_g3_6')
// (6, 7, 'lutff_4/in_3')
// (6, 7, 'sp4_h_r_46')
// (6, 7, 'sp4_r_v_b_5')
// (7, 3, 'sp4_h_r_8')
// (7, 3, 'sp4_v_t_40')
// (7, 4, 'local_g3_0')
// (7, 4, 'lutff_6/in_3')
// (7, 4, 'sp4_v_b_40')
// (7, 5, 'local_g2_5')
// (7, 5, 'lutff_6/in_3')
// (7, 5, 'sp4_v_b_29')
// (7, 6, 'sp4_h_r_5')
// (7, 6, 'sp4_v_b_16')
// (7, 7, 'local_g1_0')
// (7, 7, 'lutff_4/in_3')
// (7, 7, 'sp4_h_l_46')
// (7, 7, 'sp4_h_r_8')
// (7, 7, 'sp4_v_b_5')
// (8, 3, 'local_g1_5')
// (8, 3, 'lutff_3/in_3')
// (8, 3, 'sp4_h_r_21')
// (8, 6, 'local_g1_0')
// (8, 6, 'lutff_4/in_3')
// (8, 6, 'sp4_h_r_16')
// (8, 7, 'sp4_h_r_21')
// (9, 3, 'sp4_h_r_32')
// (9, 6, 'local_g2_5')
// (9, 6, 'lutff_4/in_3')
// (9, 6, 'sp4_h_r_29')
// (9, 7, 'sp4_h_r_32')
// (10, 3, 'sp4_h_r_45')
// (10, 3, 'sp4_r_v_b_40')
// (10, 4, 'neigh_op_tnr_0')
// (10, 4, 'sp4_r_v_b_29')
// (10, 4, 'sp4_r_v_b_45')
// (10, 5, 'neigh_op_rgt_0')
// (10, 5, 'sp4_r_v_b_16')
// (10, 5, 'sp4_r_v_b_32')
// (10, 6, 'neigh_op_bnr_0')
// (10, 6, 'sp4_h_r_40')
// (10, 6, 'sp4_r_v_b_21')
// (10, 6, 'sp4_r_v_b_5')
// (10, 7, 'sp4_h_r_45')
// (10, 7, 'sp4_r_v_b_8')
// (11, 2, 'sp4_v_t_40')
// (11, 3, 'sp4_h_l_45')
// (11, 3, 'sp4_v_b_40')
// (11, 3, 'sp4_v_t_45')
// (11, 4, 'neigh_op_top_0')
// (11, 4, 'sp4_v_b_29')
// (11, 4, 'sp4_v_b_45')
// (11, 5, 'lutff_0/out')
// (11, 5, 'sp4_v_b_16')
// (11, 5, 'sp4_v_b_32')
// (11, 6, 'neigh_op_bot_0')
// (11, 6, 'sp4_h_l_40')
// (11, 6, 'sp4_v_b_21')
// (11, 6, 'sp4_v_b_5')
// (11, 7, 'local_g1_0')
// (11, 7, 'lutff_4/in_3')
// (11, 7, 'sp4_h_l_45')
// (11, 7, 'sp4_v_b_8')
// (12, 4, 'neigh_op_tnl_0')
// (12, 5, 'neigh_op_lft_0')
// (12, 6, 'neigh_op_bnl_0')

reg n102 = 0;
// (3, 7, 'sp4_h_r_6')
// (4, 6, 'neigh_op_tnr_7')
// (4, 7, 'neigh_op_rgt_7')
// (4, 7, 'sp4_h_r_19')
// (4, 8, 'neigh_op_bnr_7')
// (5, 6, 'neigh_op_top_7')
// (5, 7, 'lutff_7/out')
// (5, 7, 'sp4_h_r_30')
// (5, 8, 'neigh_op_bot_7')
// (6, 6, 'neigh_op_tnl_7')
// (6, 7, 'local_g2_3')
// (6, 7, 'local_g3_3')
// (6, 7, 'lutff_1/in_1')
// (6, 7, 'lutff_2/in_0')
// (6, 7, 'lutff_3/in_0')
// (6, 7, 'lutff_4/in_2')
// (6, 7, 'neigh_op_lft_7')
// (6, 7, 'sp4_h_r_43')
// (6, 8, 'neigh_op_bnl_7')
// (7, 7, 'sp4_h_l_43')

wire n103;
// (3, 7, 'sp4_h_r_8')
// (4, 6, 'neigh_op_tnr_0')
// (4, 7, 'neigh_op_rgt_0')
// (4, 7, 'sp4_h_r_21')
// (4, 8, 'neigh_op_bnr_0')
// (5, 6, 'neigh_op_top_0')
// (5, 7, 'lutff_0/out')
// (5, 7, 'sp4_h_r_32')
// (5, 8, 'neigh_op_bot_0')
// (6, 6, 'neigh_op_tnl_0')
// (6, 7, 'neigh_op_lft_0')
// (6, 7, 'sp4_h_r_45')
// (6, 8, 'neigh_op_bnl_0')
// (7, 7, 'local_g0_3')
// (7, 7, 'lutff_0/in_1')
// (7, 7, 'lutff_4/in_1')
// (7, 7, 'sp4_h_l_45')
// (7, 7, 'sp4_h_r_11')
// (8, 7, 'sp4_h_r_22')
// (9, 7, 'sp4_h_r_35')
// (10, 7, 'sp4_h_r_46')
// (11, 7, 'sp4_h_l_46')

reg n104 = 0;
// (3, 7, 'sp4_r_v_b_46')
// (3, 8, 'sp4_r_v_b_35')
// (3, 9, 'sp4_r_v_b_22')
// (3, 10, 'sp4_r_v_b_11')
// (4, 6, 'sp4_h_r_5')
// (4, 6, 'sp4_v_t_46')
// (4, 7, 'sp4_v_b_46')
// (4, 8, 'sp4_v_b_35')
// (4, 9, 'sp4_v_b_22')
// (4, 10, 'local_g0_3')
// (4, 10, 'lutff_5/in_0')
// (4, 10, 'sp4_v_b_11')
// (5, 6, 'local_g1_0')
// (5, 6, 'lutff_0/in_3')
// (5, 6, 'sp4_h_r_16')
// (6, 6, 'sp12_h_r_1')
// (6, 6, 'sp4_h_r_29')
// (7, 6, 'sp12_h_r_2')
// (7, 6, 'sp4_h_r_40')
// (8, 6, 'sp12_h_r_5')
// (8, 6, 'sp4_h_l_40')
// (8, 6, 'sp4_h_r_2')
// (9, 6, 'local_g1_6')
// (9, 6, 'lutff_5/in_0')
// (9, 6, 'sp12_h_r_6')
// (9, 6, 'sp4_h_r_15')
// (10, 5, 'neigh_op_tnr_1')
// (10, 6, 'neigh_op_rgt_1')
// (10, 6, 'sp12_h_r_9')
// (10, 6, 'sp4_h_r_26')
// (10, 7, 'neigh_op_bnr_1')
// (11, 5, 'neigh_op_top_1')
// (11, 6, 'lutff_1/out')
// (11, 6, 'sp12_h_r_10')
// (11, 6, 'sp4_h_r_39')
// (11, 7, 'neigh_op_bot_1')
// (12, 5, 'neigh_op_tnl_1')
// (12, 6, 'neigh_op_lft_1')
// (12, 6, 'sp12_h_r_13')
// (12, 6, 'sp4_h_l_39')
// (12, 7, 'neigh_op_bnl_1')
// (13, 6, 'span12_horz_13')

reg n105 = 0;
// (3, 8, 'neigh_op_tnr_7')
// (3, 9, 'neigh_op_rgt_7')
// (3, 10, 'neigh_op_bnr_7')
// (4, 8, 'neigh_op_top_7')
// (4, 9, 'lutff_7/out')
// (4, 10, 'neigh_op_bot_7')
// (5, 8, 'neigh_op_tnl_7')
// (5, 9, 'local_g1_7')
// (5, 9, 'lutff_5/in_1')
// (5, 9, 'neigh_op_lft_7')
// (5, 10, 'neigh_op_bnl_7')

wire n106;
// (3, 8, 'sp4_h_r_0')
// (4, 7, 'sp4_r_v_b_43')
// (4, 8, 'local_g0_5')
// (4, 8, 'lutff_4/in_3')
// (4, 8, 'sp4_h_r_13')
// (4, 8, 'sp4_r_v_b_30')
// (4, 9, 'sp4_r_v_b_19')
// (4, 10, 'sp4_r_v_b_6')
// (5, 6, 'sp4_v_t_43')
// (5, 7, 'sp4_v_b_43')
// (5, 8, 'local_g2_0')
// (5, 8, 'lutff_5/in_3')
// (5, 8, 'lutff_7/in_3')
// (5, 8, 'sp4_h_r_24')
// (5, 8, 'sp4_v_b_30')
// (5, 9, 'local_g0_3')
// (5, 9, 'local_g1_3')
// (5, 9, 'lutff_0/in_3')
// (5, 9, 'lutff_3/in_3')
// (5, 9, 'sp4_v_b_19')
// (5, 10, 'sp4_h_r_6')
// (5, 10, 'sp4_v_b_6')
// (6, 8, 'local_g2_5')
// (6, 8, 'local_g2_6')
// (6, 8, 'lutff_1/in_3')
// (6, 8, 'lutff_2/in_3')
// (6, 8, 'sp4_h_r_37')
// (6, 8, 'sp4_r_v_b_38')
// (6, 9, 'neigh_op_tnr_7')
// (6, 9, 'sp4_r_v_b_27')
// (6, 9, 'sp4_r_v_b_43')
// (6, 10, 'neigh_op_rgt_7')
// (6, 10, 'sp4_h_r_19')
// (6, 10, 'sp4_r_v_b_14')
// (6, 10, 'sp4_r_v_b_30')
// (6, 11, 'neigh_op_bnr_7')
// (6, 11, 'sp4_r_v_b_19')
// (6, 11, 'sp4_r_v_b_3')
// (6, 12, 'sp4_r_v_b_6')
// (7, 7, 'sp4_v_t_38')
// (7, 8, 'sp4_h_l_37')
// (7, 8, 'sp4_r_v_b_39')
// (7, 8, 'sp4_v_b_38')
// (7, 8, 'sp4_v_t_43')
// (7, 9, 'neigh_op_top_7')
// (7, 9, 'sp4_r_v_b_26')
// (7, 9, 'sp4_v_b_27')
// (7, 9, 'sp4_v_b_43')
// (7, 10, 'lutff_7/out')
// (7, 10, 'sp4_h_r_30')
// (7, 10, 'sp4_r_v_b_15')
// (7, 10, 'sp4_v_b_14')
// (7, 10, 'sp4_v_b_30')
// (7, 11, 'neigh_op_bot_7')
// (7, 11, 'sp4_r_v_b_2')
// (7, 11, 'sp4_v_b_19')
// (7, 11, 'sp4_v_b_3')
// (7, 12, 'sp4_v_b_6')
// (8, 7, 'sp4_v_t_39')
// (8, 8, 'local_g2_7')
// (8, 8, 'lutff_0/in_3')
// (8, 8, 'sp4_v_b_39')
// (8, 9, 'neigh_op_tnl_7')
// (8, 9, 'sp4_v_b_26')
// (8, 10, 'neigh_op_lft_7')
// (8, 10, 'sp4_h_r_43')
// (8, 10, 'sp4_v_b_15')
// (8, 11, 'neigh_op_bnl_7')
// (8, 11, 'sp4_v_b_2')
// (9, 10, 'sp4_h_l_43')

reg n107 = 0;
// (3, 8, 'sp4_h_r_6')
// (4, 8, 'sp4_h_r_19')
// (5, 8, 'sp4_h_r_30')
// (6, 5, 'local_g2_6')
// (6, 5, 'lutff_3/in_3')
// (6, 5, 'sp4_r_v_b_37')
// (6, 5, 'sp4_r_v_b_38')
// (6, 6, 'sp4_r_v_b_24')
// (6, 6, 'sp4_r_v_b_27')
// (6, 7, 'local_g2_5')
// (6, 7, 'local_g2_6')
// (6, 7, 'lutff_1/in_3')
// (6, 7, 'lutff_2/in_3')
// (6, 7, 'lutff_3/in_2')
// (6, 7, 'sp4_r_v_b_13')
// (6, 7, 'sp4_r_v_b_14')
// (6, 8, 'sp4_h_r_43')
// (6, 8, 'sp4_r_v_b_0')
// (6, 8, 'sp4_r_v_b_3')
// (7, 3, 'local_g3_2')
// (7, 3, 'lutff_2/in_3')
// (7, 3, 'sp4_r_v_b_38')
// (7, 3, 'sp4_r_v_b_42')
// (7, 4, 'local_g0_7')
// (7, 4, 'local_g1_7')
// (7, 4, 'lutff_1/in_3')
// (7, 4, 'lutff_5/in_2')
// (7, 4, 'sp4_r_v_b_27')
// (7, 4, 'sp4_r_v_b_31')
// (7, 4, 'sp4_v_t_37')
// (7, 4, 'sp4_v_t_38')
// (7, 5, 'local_g2_6')
// (7, 5, 'lutff_1/in_3')
// (7, 5, 'lutff_2/in_2')
// (7, 5, 'sp4_r_v_b_14')
// (7, 5, 'sp4_r_v_b_18')
// (7, 5, 'sp4_r_v_b_40')
// (7, 5, 'sp4_v_b_37')
// (7, 5, 'sp4_v_b_38')
// (7, 6, 'local_g0_5')
// (7, 6, 'lutff_4/in_3')
// (7, 6, 'sp4_r_v_b_29')
// (7, 6, 'sp4_r_v_b_3')
// (7, 6, 'sp4_r_v_b_7')
// (7, 6, 'sp4_v_b_24')
// (7, 6, 'sp4_v_b_27')
// (7, 7, 'local_g2_6')
// (7, 7, 'local_g3_0')
// (7, 7, 'lutff_1/in_3')
// (7, 7, 'lutff_7/in_2')
// (7, 7, 'sp4_r_v_b_16')
// (7, 7, 'sp4_r_v_b_38')
// (7, 7, 'sp4_v_b_13')
// (7, 7, 'sp4_v_b_14')
// (7, 8, 'sp4_h_l_43')
// (7, 8, 'sp4_h_r_3')
// (7, 8, 'sp4_r_v_b_27')
// (7, 8, 'sp4_r_v_b_5')
// (7, 8, 'sp4_v_b_0')
// (7, 8, 'sp4_v_b_3')
// (7, 9, 'sp4_r_v_b_14')
// (7, 10, 'sp4_r_v_b_3')
// (8, 0, 'span12_vert_21')
// (8, 1, 'sp12_v_b_21')
// (8, 2, 'sp12_v_b_18')
// (8, 2, 'sp4_v_t_38')
// (8, 2, 'sp4_v_t_42')
// (8, 3, 'local_g3_1')
// (8, 3, 'lutff_1/in_3')
// (8, 3, 'lutff_6/in_2')
// (8, 3, 'sp12_v_b_17')
// (8, 3, 'sp4_v_b_38')
// (8, 3, 'sp4_v_b_42')
// (8, 4, 'sp12_v_b_14')
// (8, 4, 'sp4_v_b_27')
// (8, 4, 'sp4_v_b_31')
// (8, 4, 'sp4_v_t_40')
// (8, 5, 'local_g3_5')
// (8, 5, 'lutff_5/in_3')
// (8, 5, 'lutff_6/in_2')
// (8, 5, 'sp12_v_b_13')
// (8, 5, 'sp4_v_b_14')
// (8, 5, 'sp4_v_b_18')
// (8, 5, 'sp4_v_b_40')
// (8, 6, 'local_g2_2')
// (8, 6, 'lutff_1/in_3')
// (8, 6, 'sp12_v_b_10')
// (8, 6, 'sp4_h_r_8')
// (8, 6, 'sp4_v_b_29')
// (8, 6, 'sp4_v_b_3')
// (8, 6, 'sp4_v_b_7')
// (8, 6, 'sp4_v_t_38')
// (8, 7, 'sp12_v_b_9')
// (8, 7, 'sp4_v_b_16')
// (8, 7, 'sp4_v_b_38')
// (8, 8, 'sp12_v_b_6')
// (8, 8, 'sp4_h_r_14')
// (8, 8, 'sp4_v_b_27')
// (8, 8, 'sp4_v_b_5')
// (8, 9, 'sp12_v_b_5')
// (8, 9, 'sp4_v_b_14')
// (8, 10, 'sp12_v_b_2')
// (8, 10, 'sp4_v_b_3')
// (8, 11, 'sp12_h_r_1')
// (8, 11, 'sp12_v_b_1')
// (9, 3, 'local_g3_2')
// (9, 3, 'lutff_4/in_3')
// (9, 3, 'sp4_r_v_b_42')
// (9, 4, 'sp4_r_v_b_31')
// (9, 5, 'sp4_r_v_b_18')
// (9, 6, 'local_g0_5')
// (9, 6, 'lutff_0/in_3')
// (9, 6, 'lutff_3/in_2')
// (9, 6, 'lutff_6/in_3')
// (9, 6, 'sp4_h_r_21')
// (9, 6, 'sp4_r_v_b_7')
// (9, 7, 'local_g2_6')
// (9, 7, 'local_g3_2')
// (9, 7, 'lutff_1/in_3')
// (9, 7, 'lutff_3/in_3')
// (9, 7, 'lutff_5/in_2')
// (9, 7, 'sp4_r_v_b_38')
// (9, 7, 'sp4_r_v_b_42')
// (9, 8, 'sp4_h_r_27')
// (9, 8, 'sp4_r_v_b_27')
// (9, 8, 'sp4_r_v_b_31')
// (9, 9, 'sp4_r_v_b_14')
// (9, 9, 'sp4_r_v_b_18')
// (9, 10, 'sp4_r_v_b_3')
// (9, 10, 'sp4_r_v_b_7')
// (9, 11, 'sp12_h_r_2')
// (10, 2, 'sp4_h_r_7')
// (10, 2, 'sp4_v_t_42')
// (10, 3, 'sp4_v_b_42')
// (10, 4, 'sp4_v_b_31')
// (10, 5, 'sp4_v_b_18')
// (10, 6, 'sp4_h_r_32')
// (10, 6, 'sp4_v_b_7')
// (10, 6, 'sp4_v_t_38')
// (10, 6, 'sp4_v_t_42')
// (10, 7, 'sp4_v_b_38')
// (10, 7, 'sp4_v_b_42')
// (10, 8, 'sp4_h_r_38')
// (10, 8, 'sp4_v_b_27')
// (10, 8, 'sp4_v_b_31')
// (10, 9, 'sp4_r_v_b_38')
// (10, 9, 'sp4_v_b_14')
// (10, 9, 'sp4_v_b_18')
// (10, 10, 'neigh_op_tnr_7')
// (10, 10, 'sp4_r_v_b_27')
// (10, 10, 'sp4_v_b_3')
// (10, 10, 'sp4_v_b_7')
// (10, 11, 'neigh_op_rgt_7')
// (10, 11, 'sp12_h_r_5')
// (10, 11, 'sp4_r_v_b_14')
// (10, 12, 'neigh_op_bnr_7')
// (10, 12, 'sp4_r_v_b_3')
// (11, 2, 'sp4_h_r_18')
// (11, 3, 'sp4_r_v_b_39')
// (11, 4, 'sp4_r_v_b_26')
// (11, 5, 'local_g2_7')
// (11, 5, 'lutff_0/in_3')
// (11, 5, 'sp4_r_v_b_15')
// (11, 6, 'local_g2_5')
// (11, 6, 'lutff_0/in_3')
// (11, 6, 'sp4_h_r_45')
// (11, 6, 'sp4_r_v_b_2')
// (11, 8, 'sp4_h_l_38')
// (11, 8, 'sp4_v_t_38')
// (11, 9, 'sp4_v_b_38')
// (11, 10, 'neigh_op_top_7')
// (11, 10, 'sp4_v_b_27')
// (11, 11, 'lutff_7/out')
// (11, 11, 'sp12_h_r_6')
// (11, 11, 'sp4_v_b_14')
// (11, 12, 'neigh_op_bot_7')
// (11, 12, 'sp4_v_b_3')
// (12, 2, 'sp4_h_r_31')
// (12, 2, 'sp4_h_r_7')
// (12, 2, 'sp4_v_t_39')
// (12, 3, 'sp4_v_b_39')
// (12, 4, 'sp4_v_b_26')
// (12, 5, 'sp4_v_b_15')
// (12, 6, 'sp4_h_l_45')
// (12, 6, 'sp4_v_b_2')
// (12, 10, 'neigh_op_tnl_7')
// (12, 11, 'neigh_op_lft_7')
// (12, 11, 'sp12_h_r_9')
// (12, 12, 'neigh_op_bnl_7')
// (13, 2, 'span4_horz_31')
// (13, 2, 'span4_horz_7')
// (13, 11, 'span12_horz_9')

reg n108 = 0;
// (3, 8, 'sp4_r_v_b_43')
// (3, 9, 'sp4_r_v_b_30')
// (3, 10, 'neigh_op_tnr_3')
// (3, 10, 'sp4_r_v_b_19')
// (3, 11, 'neigh_op_rgt_3')
// (3, 11, 'sp4_r_v_b_6')
// (3, 12, 'neigh_op_bnr_3')
// (4, 4, 'sp4_r_v_b_42')
// (4, 5, 'sp4_r_v_b_31')
// (4, 6, 'sp4_r_v_b_18')
// (4, 7, 'sp4_r_v_b_7')
// (4, 7, 'sp4_v_t_43')
// (4, 8, 'local_g2_3')
// (4, 8, 'lutff_5/in_0')
// (4, 8, 'sp4_r_v_b_42')
// (4, 8, 'sp4_v_b_43')
// (4, 9, 'sp4_r_v_b_31')
// (4, 9, 'sp4_v_b_30')
// (4, 10, 'local_g1_3')
// (4, 10, 'lutff_2/in_0')
// (4, 10, 'neigh_op_top_3')
// (4, 10, 'sp4_r_v_b_18')
// (4, 10, 'sp4_v_b_19')
// (4, 11, 'lutff_3/out')
// (4, 11, 'sp4_r_v_b_7')
// (4, 11, 'sp4_v_b_6')
// (4, 12, 'neigh_op_bot_3')
// (5, 3, 'sp4_v_t_42')
// (5, 4, 'sp4_v_b_42')
// (5, 5, 'sp4_v_b_31')
// (5, 6, 'sp4_v_b_18')
// (5, 7, 'local_g0_7')
// (5, 7, 'lutff_0/in_3')
// (5, 7, 'sp4_v_b_7')
// (5, 7, 'sp4_v_t_42')
// (5, 8, 'sp4_v_b_42')
// (5, 9, 'sp4_v_b_31')
// (5, 10, 'neigh_op_tnl_3')
// (5, 10, 'sp4_v_b_18')
// (5, 11, 'neigh_op_lft_3')
// (5, 11, 'sp4_v_b_7')
// (5, 12, 'neigh_op_bnl_3')

reg n109 = 0;
// (3, 8, 'sp4_r_v_b_44')
// (3, 9, 'neigh_op_tnr_2')
// (3, 9, 'sp4_r_v_b_33')
// (3, 10, 'neigh_op_rgt_2')
// (3, 10, 'sp4_r_v_b_20')
// (3, 11, 'neigh_op_bnr_2')
// (3, 11, 'sp4_r_v_b_9')
// (4, 7, 'sp4_v_t_44')
// (4, 8, 'sp4_v_b_44')
// (4, 9, 'neigh_op_top_2')
// (4, 9, 'sp4_v_b_33')
// (4, 10, 'lutff_2/out')
// (4, 10, 'sp4_v_b_20')
// (4, 11, 'local_g0_1')
// (4, 11, 'lutff_0/in_1')
// (4, 11, 'neigh_op_bot_2')
// (4, 11, 'sp4_v_b_9')
// (5, 9, 'neigh_op_tnl_2')
// (5, 10, 'neigh_op_lft_2')
// (5, 11, 'neigh_op_bnl_2')

reg n110 = 0;
// (3, 9, 'neigh_op_tnr_3')
// (3, 10, 'neigh_op_rgt_3')
// (3, 11, 'neigh_op_bnr_3')
// (4, 9, 'neigh_op_top_3')
// (4, 10, 'lutff_3/out')
// (4, 11, 'neigh_op_bot_3')
// (5, 9, 'neigh_op_tnl_3')
// (5, 10, 'neigh_op_lft_3')
// (5, 11, 'local_g2_3')
// (5, 11, 'lutff_0/in_3')
// (5, 11, 'neigh_op_bnl_3')

reg n111 = 0;
// (3, 9, 'neigh_op_tnr_6')
// (3, 10, 'neigh_op_rgt_6')
// (3, 11, 'neigh_op_bnr_6')
// (4, 9, 'neigh_op_top_6')
// (4, 10, 'lutff_6/out')
// (4, 11, 'neigh_op_bot_6')
// (5, 9, 'neigh_op_tnl_6')
// (5, 10, 'neigh_op_lft_6')
// (5, 11, 'local_g2_6')
// (5, 11, 'lutff_3/in_3')
// (5, 11, 'neigh_op_bnl_6')

wire n112;
// (3, 9, 'sp4_h_r_10')
// (4, 8, 'neigh_op_tnr_1')
// (4, 9, 'neigh_op_rgt_1')
// (4, 9, 'sp4_h_r_23')
// (4, 10, 'neigh_op_bnr_1')
// (5, 8, 'neigh_op_top_1')
// (5, 9, 'lutff_1/out')
// (5, 9, 'sp4_h_r_34')
// (5, 10, 'neigh_op_bot_1')
// (6, 2, 'sp4_r_v_b_42')
// (6, 3, 'sp4_r_v_b_31')
// (6, 4, 'sp4_r_v_b_18')
// (6, 5, 'sp4_r_v_b_7')
// (6, 6, 'sp4_r_v_b_41')
// (6, 7, 'sp4_r_v_b_28')
// (6, 8, 'neigh_op_tnl_1')
// (6, 8, 'sp4_r_v_b_17')
// (6, 9, 'neigh_op_lft_1')
// (6, 9, 'sp4_h_r_47')
// (6, 9, 'sp4_r_v_b_4')
// (6, 10, 'neigh_op_bnl_1')
// (7, 1, 'sp4_v_t_42')
// (7, 2, 'sp4_v_b_42')
// (7, 3, 'sp4_v_b_31')
// (7, 4, 'local_g0_2')
// (7, 4, 'local_g1_2')
// (7, 4, 'lutff_0/in_0')
// (7, 4, 'lutff_6/in_1')
// (7, 4, 'sp4_v_b_18')
// (7, 5, 'sp4_v_b_7')
// (7, 5, 'sp4_v_t_41')
// (7, 6, 'sp4_v_b_41')
// (7, 7, 'sp4_v_b_28')
// (7, 8, 'sp4_v_b_17')
// (7, 9, 'sp4_h_l_47')
// (7, 9, 'sp4_v_b_4')

wire n113;
// (3, 10, 'neigh_op_tnr_0')
// (3, 11, 'neigh_op_rgt_0')
// (3, 12, 'neigh_op_bnr_0')
// (4, 10, 'neigh_op_top_0')
// (4, 10, 'sp4_r_v_b_44')
// (4, 11, 'lutff_0/out')
// (4, 11, 'sp4_r_v_b_33')
// (4, 12, 'neigh_op_bot_0')
// (4, 12, 'sp4_r_v_b_20')
// (4, 13, 'sp4_r_v_b_9')
// (5, 9, 'sp4_v_t_44')
// (5, 10, 'neigh_op_tnl_0')
// (5, 10, 'sp4_v_b_44')
// (5, 11, 'neigh_op_lft_0')
// (5, 11, 'sp4_v_b_33')
// (5, 12, 'neigh_op_bnl_0')
// (5, 12, 'sp4_v_b_20')
// (5, 13, 'sp4_h_r_9')
// (5, 13, 'sp4_v_b_9')
// (6, 13, 'local_g0_4')
// (6, 13, 'lutff_3/in_3')
// (6, 13, 'lutff_7/in_3')
// (6, 13, 'sp4_h_r_20')
// (7, 13, 'sp4_h_r_33')
// (8, 13, 'sp4_h_r_44')
// (9, 13, 'sp4_h_l_44')

wire n114;
// (3, 10, 'neigh_op_tnr_2')
// (3, 11, 'neigh_op_rgt_2')
// (3, 12, 'neigh_op_bnr_2')
// (4, 10, 'neigh_op_top_2')
// (4, 11, 'local_g1_2')
// (4, 11, 'lutff_0/in_3')
// (4, 11, 'lutff_2/out')
// (4, 12, 'neigh_op_bot_2')
// (5, 10, 'neigh_op_tnl_2')
// (5, 11, 'neigh_op_lft_2')
// (5, 12, 'neigh_op_bnl_2')

reg n115 = 0;
// (3, 10, 'neigh_op_tnr_6')
// (3, 11, 'neigh_op_rgt_6')
// (3, 12, 'neigh_op_bnr_6')
// (4, 10, 'neigh_op_top_6')
// (4, 11, 'local_g0_6')
// (4, 11, 'lutff_4/in_0')
// (4, 11, 'lutff_6/out')
// (4, 12, 'neigh_op_bot_6')
// (5, 10, 'neigh_op_tnl_6')
// (5, 11, 'neigh_op_lft_6')
// (5, 12, 'neigh_op_bnl_6')

wire n116;
// (3, 11, 'neigh_op_tnr_1')
// (3, 12, 'neigh_op_rgt_1')
// (3, 13, 'neigh_op_bnr_1')
// (4, 11, 'neigh_op_top_1')
// (4, 12, 'local_g0_1')
// (4, 12, 'local_g1_1')
// (4, 12, 'lutff_1/out')
// (4, 12, 'lutff_4/in_2')
// (4, 12, 'lutff_5/in_0')
// (4, 13, 'neigh_op_bot_1')
// (5, 11, 'neigh_op_tnl_1')
// (5, 12, 'neigh_op_lft_1')
// (5, 13, 'neigh_op_bnl_1')

wire n117;
// (3, 11, 'neigh_op_tnr_2')
// (3, 12, 'neigh_op_rgt_2')
// (3, 13, 'neigh_op_bnr_2')
// (4, 11, 'neigh_op_top_2')
// (4, 12, 'local_g0_2')
// (4, 12, 'local_g1_2')
// (4, 12, 'lutff_2/out')
// (4, 12, 'lutff_4/in_3')
// (4, 12, 'lutff_5/in_3')
// (4, 13, 'neigh_op_bot_2')
// (5, 11, 'neigh_op_tnl_2')
// (5, 12, 'neigh_op_lft_2')
// (5, 13, 'neigh_op_bnl_2')

wire n118;
// (3, 11, 'neigh_op_tnr_3')
// (3, 12, 'neigh_op_rgt_3')
// (3, 13, 'neigh_op_bnr_3')
// (4, 11, 'neigh_op_top_3')
// (4, 12, 'local_g0_3')
// (4, 12, 'lutff_3/out')
// (4, 12, 'lutff_5/in_2')
// (4, 13, 'neigh_op_bot_3')
// (5, 11, 'neigh_op_tnl_3')
// (5, 12, 'neigh_op_lft_3')
// (5, 13, 'neigh_op_bnl_3')

reg n119 = 0;
// (3, 11, 'neigh_op_tnr_6')
// (3, 12, 'neigh_op_rgt_6')
// (3, 13, 'neigh_op_bnr_6')
// (4, 11, 'neigh_op_top_6')
// (4, 12, 'local_g1_6')
// (4, 12, 'lutff_2/in_3')
// (4, 12, 'lutff_6/out')
// (4, 13, 'neigh_op_bot_6')
// (5, 11, 'neigh_op_tnl_6')
// (5, 12, 'neigh_op_lft_6')
// (5, 13, 'neigh_op_bnl_6')

reg n120 = 0;
// (3, 11, 'neigh_op_tnr_7')
// (3, 12, 'neigh_op_rgt_7')
// (3, 13, 'neigh_op_bnr_7')
// (4, 11, 'neigh_op_top_7')
// (4, 12, 'local_g1_7')
// (4, 12, 'lutff_3/in_3')
// (4, 12, 'lutff_7/out')
// (4, 13, 'neigh_op_bot_7')
// (5, 11, 'neigh_op_tnl_7')
// (5, 12, 'neigh_op_lft_7')
// (5, 13, 'neigh_op_bnl_7')

wire n121;
// (3, 11, 'sp4_r_v_b_38')
// (3, 12, 'neigh_op_tnr_7')
// (3, 12, 'sp4_r_v_b_27')
// (3, 13, 'neigh_op_rgt_7')
// (3, 13, 'sp4_r_v_b_14')
// (3, 14, 'neigh_op_bnr_7')
// (3, 14, 'sp4_r_v_b_3')
// (4, 10, 'sp4_v_t_38')
// (4, 11, 'sp4_v_b_38')
// (4, 12, 'neigh_op_top_7')
// (4, 12, 'sp4_v_b_27')
// (4, 13, 'lutff_7/out')
// (4, 13, 'sp4_v_b_14')
// (4, 14, 'local_g1_3')
// (4, 14, 'lutff_global/cen')
// (4, 14, 'neigh_op_bot_7')
// (4, 14, 'sp4_v_b_3')
// (5, 12, 'neigh_op_tnl_7')
// (5, 13, 'neigh_op_lft_7')
// (5, 14, 'neigh_op_bnl_7')

wire n122;
// (3, 12, 'sp4_h_r_7')
// (4, 12, 'sp4_h_r_18')
// (5, 11, 'neigh_op_tnr_5')
// (5, 12, 'neigh_op_rgt_5')
// (5, 12, 'sp4_h_r_31')
// (5, 13, 'neigh_op_bnr_5')
// (6, 11, 'neigh_op_top_5')
// (6, 12, 'lutff_5/out')
// (6, 12, 'sp4_h_r_42')
// (6, 13, 'local_g0_5')
// (6, 13, 'lutff_4/in_1')
// (6, 13, 'lutff_6/in_3')
// (6, 13, 'neigh_op_bot_5')
// (6, 13, 'sp4_r_v_b_42')
// (6, 14, 'sp4_r_v_b_31')
// (6, 15, 'sp4_r_v_b_18')
// (6, 16, 'sp4_r_v_b_7')
// (7, 11, 'neigh_op_tnl_5')
// (7, 12, 'neigh_op_lft_5')
// (7, 12, 'sp4_h_l_42')
// (7, 12, 'sp4_v_t_42')
// (7, 13, 'local_g3_2')
// (7, 13, 'local_g3_5')
// (7, 13, 'lutff_1/in_3')
// (7, 13, 'lutff_4/in_1')
// (7, 13, 'neigh_op_bnl_5')
// (7, 13, 'sp4_v_b_42')
// (7, 14, 'sp4_v_b_31')
// (7, 15, 'sp4_v_b_18')
// (7, 16, 'sp4_v_b_7')

reg n123 = 0;
// (3, 12, 'sp4_r_v_b_36')
// (3, 13, 'sp4_r_v_b_25')
// (3, 14, 'sp4_r_v_b_12')
// (3, 15, 'sp4_r_v_b_1')
// (4, 2, 'sp12_v_t_22')
// (4, 3, 'sp12_v_b_22')
// (4, 4, 'sp12_v_b_21')
// (4, 5, 'sp12_v_b_18')
// (4, 6, 'sp12_v_b_17')
// (4, 7, 'sp12_v_b_14')
// (4, 8, 'sp12_v_b_13')
// (4, 9, 'sp12_v_b_10')
// (4, 10, 'sp12_v_b_9')
// (4, 11, 'sp12_v_b_6')
// (4, 11, 'sp4_v_t_36')
// (4, 12, 'sp12_v_b_5')
// (4, 12, 'sp4_v_b_36')
// (4, 13, 'local_g3_2')
// (4, 13, 'lutff_7/in_2')
// (4, 13, 'sp12_v_b_2')
// (4, 13, 'sp4_v_b_25')
// (4, 14, 'local_g1_1')
// (4, 14, 'lutff_5/in_1')
// (4, 14, 'sp12_h_r_1')
// (4, 14, 'sp12_v_b_1')
// (4, 14, 'sp4_v_b_12')
// (4, 15, 'local_g0_1')
// (4, 15, 'local_g1_1')
// (4, 15, 'lutff_3/in_0')
// (4, 15, 'lutff_7/in_1')
// (4, 15, 'sp4_v_b_1')
// (5, 14, 'sp12_h_r_2')
// (6, 14, 'sp12_h_r_5')
// (7, 14, 'sp12_h_r_6')
// (8, 13, 'neigh_op_tnr_1')
// (8, 14, 'neigh_op_rgt_1')
// (8, 14, 'sp12_h_r_9')
// (8, 15, 'neigh_op_bnr_1')
// (9, 11, 'sp12_h_r_1')
// (9, 11, 'sp12_v_t_22')
// (9, 12, 'sp12_v_b_22')
// (9, 13, 'neigh_op_top_1')
// (9, 13, 'sp12_v_b_21')
// (9, 14, 'local_g0_1')
// (9, 14, 'lutff_1/in_2')
// (9, 14, 'lutff_1/out')
// (9, 14, 'sp12_h_r_10')
// (9, 14, 'sp12_v_b_18')
// (9, 15, 'neigh_op_bot_1')
// (9, 15, 'sp12_v_b_17')
// (9, 16, 'sp12_v_b_14')
// (9, 17, 'span12_vert_13')
// (10, 11, 'sp12_h_r_2')
// (10, 13, 'neigh_op_tnl_1')
// (10, 14, 'neigh_op_lft_1')
// (10, 14, 'sp12_h_r_13')
// (10, 15, 'neigh_op_bnl_1')
// (11, 11, 'local_g1_5')
// (11, 11, 'lutff_global/s_r')
// (11, 11, 'sp12_h_r_5')
// (11, 14, 'sp12_h_r_14')
// (12, 11, 'sp12_h_r_6')
// (12, 14, 'sp12_h_r_17')
// (13, 11, 'span12_horz_6')
// (13, 14, 'span12_horz_17')

reg n124 = 0;
// (3, 13, 'neigh_op_tnr_2')
// (3, 14, 'neigh_op_rgt_2')
// (3, 15, 'neigh_op_bnr_2')
// (4, 13, 'neigh_op_top_2')
// (4, 14, 'local_g0_2')
// (4, 14, 'lutff_2/in_2')
// (4, 14, 'lutff_2/out')
// (4, 15, 'local_g0_2')
// (4, 15, 'local_g1_2')
// (4, 15, 'lutff_1/in_0')
// (4, 15, 'lutff_2/in_0')
// (4, 15, 'lutff_4/in_1')
// (4, 15, 'lutff_6/in_0')
// (4, 15, 'neigh_op_bot_2')
// (5, 13, 'neigh_op_tnl_2')
// (5, 14, 'neigh_op_lft_2')
// (5, 15, 'neigh_op_bnl_2')

reg n125 = 0;
// (3, 13, 'neigh_op_tnr_3')
// (3, 14, 'neigh_op_rgt_3')
// (3, 15, 'neigh_op_bnr_3')
// (4, 13, 'neigh_op_top_3')
// (4, 14, 'local_g0_3')
// (4, 14, 'lutff_3/in_2')
// (4, 14, 'lutff_3/out')
// (4, 15, 'local_g0_3')
// (4, 15, 'local_g1_3')
// (4, 15, 'lutff_1/in_1')
// (4, 15, 'lutff_2/in_1')
// (4, 15, 'lutff_4/in_0')
// (4, 15, 'lutff_6/in_1')
// (4, 15, 'neigh_op_bot_3')
// (5, 13, 'neigh_op_tnl_3')
// (5, 14, 'neigh_op_lft_3')
// (5, 15, 'neigh_op_bnl_3')

reg n126 = 0;
// (3, 13, 'neigh_op_tnr_4')
// (3, 14, 'neigh_op_rgt_4')
// (3, 15, 'neigh_op_bnr_4')
// (4, 13, 'neigh_op_top_4')
// (4, 14, 'local_g0_4')
// (4, 14, 'local_g1_4')
// (4, 14, 'lutff_1/in_2')
// (4, 14, 'lutff_4/in_2')
// (4, 14, 'lutff_4/out')
// (4, 15, 'local_g0_4')
// (4, 15, 'local_g1_4')
// (4, 15, 'lutff_1/in_2')
// (4, 15, 'lutff_2/in_2')
// (4, 15, 'lutff_4/in_2')
// (4, 15, 'lutff_6/in_2')
// (4, 15, 'neigh_op_bot_4')
// (5, 13, 'neigh_op_tnl_4')
// (5, 14, 'neigh_op_lft_4')
// (5, 15, 'neigh_op_bnl_4')

reg n127 = 0;
// (3, 13, 'neigh_op_tnr_5')
// (3, 14, 'neigh_op_rgt_5')
// (3, 15, 'neigh_op_bnr_5')
// (4, 13, 'neigh_op_top_5')
// (4, 14, 'local_g0_5')
// (4, 14, 'local_g1_5')
// (4, 14, 'lutff_0/in_1')
// (4, 14, 'lutff_4/in_3')
// (4, 14, 'lutff_5/in_3')
// (4, 14, 'lutff_5/out')
// (4, 15, 'local_g0_5')
// (4, 15, 'local_g1_5')
// (4, 15, 'lutff_1/in_3')
// (4, 15, 'lutff_2/in_3')
// (4, 15, 'lutff_4/in_3')
// (4, 15, 'lutff_6/in_3')
// (4, 15, 'neigh_op_bot_5')
// (5, 13, 'neigh_op_tnl_5')
// (5, 14, 'neigh_op_lft_5')
// (5, 15, 'neigh_op_bnl_5')

wire n128;
// (3, 14, 'neigh_op_tnr_0')
// (3, 15, 'neigh_op_rgt_0')
// (3, 16, 'neigh_op_bnr_0')
// (4, 14, 'neigh_op_top_0')
// (4, 15, 'local_g2_0')
// (4, 15, 'lutff_0/out')
// (4, 15, 'lutff_3/in_3')
// (4, 16, 'neigh_op_bot_0')
// (5, 14, 'neigh_op_tnl_0')
// (5, 15, 'neigh_op_lft_0')
// (5, 16, 'neigh_op_bnl_0')

wire n129;
// (3, 14, 'neigh_op_tnr_2')
// (3, 15, 'neigh_op_rgt_2')
// (3, 16, 'neigh_op_bnr_2')
// (4, 13, 'sp4_r_v_b_45')
// (4, 14, 'neigh_op_top_2')
// (4, 14, 'sp4_r_v_b_32')
// (4, 15, 'local_g3_5')
// (4, 15, 'lutff_0/in_0')
// (4, 15, 'lutff_2/out')
// (4, 15, 'sp4_r_v_b_21')
// (4, 16, 'neigh_op_bot_2')
// (4, 16, 'sp4_r_v_b_8')
// (5, 12, 'sp4_v_t_45')
// (5, 13, 'sp4_v_b_45')
// (5, 14, 'neigh_op_tnl_2')
// (5, 14, 'sp4_v_b_32')
// (5, 15, 'local_g0_2')
// (5, 15, 'local_g1_2')
// (5, 15, 'lutff_0/in_2')
// (5, 15, 'lutff_7/in_0')
// (5, 15, 'neigh_op_lft_2')
// (5, 15, 'sp4_v_b_21')
// (5, 16, 'neigh_op_bnl_2')
// (5, 16, 'sp4_v_b_8')

wire n130;
// (3, 14, 'neigh_op_tnr_3')
// (3, 15, 'neigh_op_rgt_3')
// (3, 16, 'neigh_op_bnr_3')
// (4, 13, 'sp4_r_v_b_47')
// (4, 14, 'local_g0_1')
// (4, 14, 'local_g2_2')
// (4, 14, 'lutff_2/in_0')
// (4, 14, 'lutff_3/in_0')
// (4, 14, 'lutff_4/in_0')
// (4, 14, 'neigh_op_top_3')
// (4, 14, 'sp4_r_v_b_34')
// (4, 15, 'lutff_3/out')
// (4, 15, 'sp4_r_v_b_23')
// (4, 16, 'neigh_op_bot_3')
// (4, 16, 'sp4_r_v_b_10')
// (5, 12, 'sp4_v_t_47')
// (5, 13, 'sp4_v_b_47')
// (5, 14, 'neigh_op_tnl_3')
// (5, 14, 'sp4_v_b_34')
// (5, 15, 'neigh_op_lft_3')
// (5, 15, 'sp4_v_b_23')
// (5, 16, 'neigh_op_bnl_3')
// (5, 16, 'sp4_v_b_10')

wire n131;
// (3, 14, 'neigh_op_tnr_6')
// (3, 15, 'neigh_op_rgt_6')
// (3, 16, 'neigh_op_bnr_6')
// (4, 14, 'neigh_op_top_6')
// (4, 15, 'local_g1_6')
// (4, 15, 'lutff_5/in_2')
// (4, 15, 'lutff_6/out')
// (4, 15, 'lutff_7/in_2')
// (4, 16, 'neigh_op_bot_6')
// (5, 14, 'neigh_op_tnl_6')
// (5, 15, 'neigh_op_lft_6')
// (5, 16, 'neigh_op_bnl_6')

wire n132;
// (3, 14, 'sp12_h_r_1')
// (4, 14, 'sp12_h_r_2')
// (5, 13, 'neigh_op_tnr_7')
// (5, 14, 'neigh_op_rgt_7')
// (5, 14, 'sp12_h_r_5')
// (5, 14, 'sp4_h_r_3')
// (5, 15, 'neigh_op_bnr_7')
// (6, 13, 'neigh_op_top_7')
// (6, 14, 'lutff_7/out')
// (6, 14, 'sp12_h_r_6')
// (6, 14, 'sp4_h_r_14')
// (6, 15, 'local_g1_7')
// (6, 15, 'lutff_2/in_0')
// (6, 15, 'neigh_op_bot_7')
// (7, 13, 'neigh_op_tnl_7')
// (7, 14, 'local_g0_1')
// (7, 14, 'local_g1_1')
// (7, 14, 'local_g1_4')
// (7, 14, 'lutff_1/in_0')
// (7, 14, 'lutff_2/in_3')
// (7, 14, 'lutff_6/in_2')
// (7, 14, 'lutff_7/in_2')
// (7, 14, 'neigh_op_lft_7')
// (7, 14, 'sp12_h_r_9')
// (7, 14, 'sp4_h_r_27')
// (7, 14, 'sp4_h_r_4')
// (7, 15, 'local_g3_7')
// (7, 15, 'lutff_6/in_0')
// (7, 15, 'neigh_op_bnl_7')
// (8, 14, 'local_g2_6')
// (8, 14, 'local_g3_6')
// (8, 14, 'lutff_0/in_0')
// (8, 14, 'lutff_1/in_1')
// (8, 14, 'lutff_2/in_1')
// (8, 14, 'sp12_h_r_10')
// (8, 14, 'sp4_h_r_17')
// (8, 14, 'sp4_h_r_38')
// (9, 14, 'sp12_h_r_13')
// (9, 14, 'sp4_h_l_38')
// (9, 14, 'sp4_h_r_28')
// (10, 14, 'sp12_h_r_14')
// (10, 14, 'sp4_h_r_41')
// (11, 14, 'sp12_h_r_17')
// (11, 14, 'sp4_h_l_41')
// (12, 14, 'sp12_h_r_18')
// (13, 14, 'span12_horz_18')

wire n133;
// (3, 14, 'sp4_h_r_5')
// (4, 14, 'sp4_h_r_16')
// (5, 11, 'neigh_op_tnr_6')
// (5, 12, 'neigh_op_rgt_6')
// (5, 13, 'neigh_op_bnr_6')
// (5, 14, 'sp4_h_r_29')
// (6, 11, 'neigh_op_top_6')
// (6, 11, 'sp4_r_v_b_40')
// (6, 12, 'lutff_6/out')
// (6, 12, 'sp4_r_v_b_29')
// (6, 13, 'neigh_op_bot_6')
// (6, 13, 'sp4_r_v_b_16')
// (6, 14, 'local_g1_5')
// (6, 14, 'lutff_0/in_2')
// (6, 14, 'lutff_4/in_2')
// (6, 14, 'sp4_h_r_40')
// (6, 14, 'sp4_r_v_b_5')
// (7, 10, 'sp4_v_t_40')
// (7, 11, 'neigh_op_tnl_6')
// (7, 11, 'sp4_v_b_40')
// (7, 12, 'neigh_op_lft_6')
// (7, 12, 'sp4_v_b_29')
// (7, 13, 'local_g3_6')
// (7, 13, 'lutff_2/in_3')
// (7, 13, 'neigh_op_bnl_6')
// (7, 13, 'sp4_v_b_16')
// (7, 14, 'local_g0_0')
// (7, 14, 'lutff_4/in_2')
// (7, 14, 'sp4_h_l_40')
// (7, 14, 'sp4_h_r_8')
// (7, 14, 'sp4_v_b_5')
// (8, 14, 'sp4_h_r_21')
// (9, 14, 'sp4_h_r_32')
// (10, 14, 'sp4_h_r_45')
// (11, 14, 'sp4_h_l_45')

reg \d_out[5] = 0 ;
// (4, 1, 'sp4_r_v_b_45')
// (4, 2, 'sp4_r_v_b_32')
// (4, 3, 'neigh_op_tnr_4')
// (4, 3, 'sp4_r_v_b_21')
// (4, 4, 'neigh_op_rgt_4')
// (4, 4, 'sp4_r_v_b_8')
// (4, 5, 'neigh_op_bnr_4')
// (5, 0, 'io_0/D_OUT_0')
// (5, 0, 'io_0/PAD')
// (5, 0, 'local_g1_5')
// (5, 0, 'span4_vert_45')
// (5, 1, 'sp4_v_b_45')
// (5, 2, 'sp4_v_b_32')
// (5, 3, 'neigh_op_top_4')
// (5, 3, 'sp4_v_b_21')
// (5, 4, 'lutff_4/out')
// (5, 4, 'sp4_v_b_8')
// (5, 5, 'neigh_op_bot_4')
// (6, 3, 'neigh_op_tnl_4')
// (6, 4, 'neigh_op_lft_4')
// (6, 5, 'neigh_op_bnl_4')

reg n135 = 0;
// (4, 2, 'neigh_op_tnr_1')
// (4, 3, 'neigh_op_rgt_1')
// (4, 4, 'neigh_op_bnr_1')
// (5, 2, 'neigh_op_top_1')
// (5, 3, 'local_g1_1')
// (5, 3, 'lutff_1/out')
// (5, 3, 'lutff_2/in_0')
// (5, 4, 'neigh_op_bot_1')
// (6, 2, 'neigh_op_tnl_1')
// (6, 3, 'neigh_op_lft_1')
// (6, 4, 'neigh_op_bnl_1')

reg n136 = 0;
// (4, 2, 'neigh_op_tnr_2')
// (4, 3, 'neigh_op_rgt_2')
// (4, 4, 'neigh_op_bnr_2')
// (5, 2, 'neigh_op_top_2')
// (5, 3, 'local_g1_2')
// (5, 3, 'lutff_2/out')
// (5, 3, 'lutff_7/in_0')
// (5, 4, 'neigh_op_bot_2')
// (6, 2, 'neigh_op_tnl_2')
// (6, 3, 'neigh_op_lft_2')
// (6, 4, 'neigh_op_bnl_2')

reg n137 = 0;
// (4, 2, 'neigh_op_tnr_3')
// (4, 3, 'local_g3_3')
// (4, 3, 'lutff_4/in_0')
// (4, 3, 'neigh_op_rgt_3')
// (4, 4, 'neigh_op_bnr_3')
// (5, 2, 'neigh_op_top_3')
// (5, 3, 'lutff_3/out')
// (5, 4, 'neigh_op_bot_3')
// (6, 2, 'neigh_op_tnl_3')
// (6, 3, 'neigh_op_lft_3')
// (6, 4, 'neigh_op_bnl_3')

reg n138 = 0;
// (4, 2, 'neigh_op_tnr_5')
// (4, 3, 'neigh_op_rgt_5')
// (4, 4, 'neigh_op_bnr_5')
// (5, 2, 'neigh_op_top_5')
// (5, 3, 'local_g0_5')
// (5, 3, 'lutff_3/in_0')
// (5, 3, 'lutff_5/out')
// (5, 4, 'neigh_op_bot_5')
// (6, 2, 'neigh_op_tnl_5')
// (6, 3, 'neigh_op_lft_5')
// (6, 4, 'neigh_op_bnl_5')

reg n139 = 0;
// (4, 2, 'neigh_op_tnr_6')
// (4, 3, 'neigh_op_rgt_6')
// (4, 4, 'neigh_op_bnr_6')
// (5, 2, 'neigh_op_top_6')
// (5, 3, 'lutff_6/out')
// (5, 4, 'local_g1_6')
// (5, 4, 'lutff_2/in_3')
// (5, 4, 'neigh_op_bot_6')
// (6, 2, 'neigh_op_tnl_6')
// (6, 3, 'neigh_op_lft_6')
// (6, 4, 'neigh_op_bnl_6')

reg n140 = 0;
// (4, 2, 'neigh_op_tnr_7')
// (4, 3, 'neigh_op_rgt_7')
// (4, 4, 'neigh_op_bnr_7')
// (5, 2, 'neigh_op_top_7')
// (5, 3, 'local_g1_7')
// (5, 3, 'lutff_6/in_0')
// (5, 3, 'lutff_7/out')
// (5, 4, 'neigh_op_bot_7')
// (6, 2, 'neigh_op_tnl_7')
// (6, 3, 'neigh_op_lft_7')
// (6, 4, 'neigh_op_bnl_7')

reg n141 = 0;
// (4, 3, 'neigh_op_tnr_0')
// (4, 4, 'neigh_op_rgt_0')
// (4, 5, 'neigh_op_bnr_0')
// (5, 3, 'neigh_op_top_0')
// (5, 4, 'local_g1_0')
// (5, 4, 'lutff_0/out')
// (5, 4, 'lutff_1/in_0')
// (5, 5, 'neigh_op_bot_0')
// (6, 3, 'neigh_op_tnl_0')
// (6, 4, 'neigh_op_lft_0')
// (6, 5, 'neigh_op_bnl_0')

reg n142 = 0;
// (4, 3, 'neigh_op_tnr_2')
// (4, 4, 'neigh_op_rgt_2')
// (4, 5, 'neigh_op_bnr_2')
// (5, 3, 'neigh_op_top_2')
// (5, 4, 'lutff_2/out')
// (5, 4, 'sp4_h_r_4')
// (5, 5, 'neigh_op_bot_2')
// (6, 3, 'neigh_op_tnl_2')
// (6, 4, 'local_g1_1')
// (6, 4, 'lutff_2/in_0')
// (6, 4, 'neigh_op_lft_2')
// (6, 4, 'sp4_h_r_17')
// (6, 5, 'neigh_op_bnl_2')
// (7, 4, 'sp4_h_r_28')
// (8, 4, 'sp4_h_r_41')
// (9, 4, 'sp4_h_l_41')

reg n143 = 0;
// (4, 3, 'neigh_op_tnr_3')
// (4, 4, 'neigh_op_rgt_3')
// (4, 5, 'neigh_op_bnr_3')
// (5, 1, 'sp4_r_v_b_42')
// (5, 2, 'sp4_r_v_b_31')
// (5, 3, 'neigh_op_top_3')
// (5, 3, 'sp4_r_v_b_18')
// (5, 4, 'lutff_3/out')
// (5, 4, 'sp4_r_v_b_7')
// (5, 5, 'neigh_op_bot_3')
// (6, 0, 'span4_vert_42')
// (6, 1, 'sp4_v_b_42')
// (6, 2, 'sp4_v_b_31')
// (6, 3, 'neigh_op_tnl_3')
// (6, 3, 'sp4_v_b_18')
// (6, 4, 'local_g1_7')
// (6, 4, 'lutff_0/in_0')
// (6, 4, 'neigh_op_lft_3')
// (6, 4, 'sp4_v_b_7')
// (6, 5, 'neigh_op_bnl_3')

reg n144 = 0;
// (4, 3, 'neigh_op_tnr_5')
// (4, 4, 'neigh_op_rgt_5')
// (4, 5, 'neigh_op_bnr_5')
// (5, 3, 'neigh_op_top_5')
// (5, 4, 'local_g0_5')
// (5, 4, 'lutff_5/out')
// (5, 4, 'lutff_7/in_0')
// (5, 5, 'neigh_op_bot_5')
// (6, 3, 'neigh_op_tnl_5')
// (6, 4, 'neigh_op_lft_5')
// (6, 5, 'neigh_op_bnl_5')

reg n145 = 0;
// (4, 3, 'neigh_op_tnr_6')
// (4, 4, 'neigh_op_rgt_6')
// (4, 5, 'neigh_op_bnr_6')
// (5, 3, 'neigh_op_top_6')
// (5, 4, 'local_g3_6')
// (5, 4, 'lutff_0/in_3')
// (5, 4, 'lutff_6/out')
// (5, 5, 'neigh_op_bot_6')
// (6, 3, 'neigh_op_tnl_6')
// (6, 4, 'neigh_op_lft_6')
// (6, 5, 'neigh_op_bnl_6')

reg n146 = 0;
// (4, 3, 'neigh_op_tnr_7')
// (4, 4, 'local_g3_7')
// (4, 4, 'lutff_1/in_3')
// (4, 4, 'neigh_op_rgt_7')
// (4, 5, 'neigh_op_bnr_7')
// (5, 3, 'neigh_op_top_7')
// (5, 4, 'local_g0_7')
// (5, 4, 'local_g1_7')
// (5, 4, 'lutff_0/in_2')
// (5, 4, 'lutff_4/in_3')
// (5, 4, 'lutff_7/out')
// (5, 5, 'neigh_op_bot_7')
// (6, 3, 'neigh_op_tnl_7')
// (6, 4, 'neigh_op_lft_7')
// (6, 5, 'neigh_op_bnl_7')

reg n147 = 0;
// (4, 4, 'neigh_op_tnr_0')
// (4, 5, 'neigh_op_rgt_0')
// (4, 6, 'neigh_op_bnr_0')
// (5, 4, 'neigh_op_top_0')
// (5, 5, 'local_g1_0')
// (5, 5, 'lutff_0/out')
// (5, 5, 'lutff_7/in_0')
// (5, 6, 'neigh_op_bot_0')
// (6, 4, 'neigh_op_tnl_0')
// (6, 5, 'neigh_op_lft_0')
// (6, 6, 'neigh_op_bnl_0')

reg n148 = 0;
// (4, 4, 'neigh_op_tnr_1')
// (4, 5, 'neigh_op_rgt_1')
// (4, 6, 'neigh_op_bnr_1')
// (5, 4, 'neigh_op_top_1')
// (5, 5, 'local_g0_1')
// (5, 5, 'lutff_1/out')
// (5, 5, 'lutff_5/in_0')
// (5, 6, 'neigh_op_bot_1')
// (6, 4, 'neigh_op_tnl_1')
// (6, 5, 'neigh_op_lft_1')
// (6, 6, 'neigh_op_bnl_1')

reg n149 = 0;
// (4, 4, 'neigh_op_tnr_2')
// (4, 5, 'neigh_op_rgt_2')
// (4, 6, 'neigh_op_bnr_2')
// (5, 4, 'neigh_op_top_2')
// (5, 5, 'local_g0_2')
// (5, 5, 'lutff_2/out')
// (5, 5, 'lutff_6/in_0')
// (5, 6, 'neigh_op_bot_2')
// (6, 4, 'neigh_op_tnl_2')
// (6, 5, 'neigh_op_lft_2')
// (6, 6, 'neigh_op_bnl_2')

reg n150 = 0;
// (4, 4, 'neigh_op_tnr_3')
// (4, 5, 'neigh_op_rgt_3')
// (4, 6, 'neigh_op_bnr_3')
// (5, 4, 'neigh_op_top_3')
// (5, 5, 'local_g0_3')
// (5, 5, 'lutff_1/in_0')
// (5, 5, 'lutff_3/out')
// (5, 6, 'neigh_op_bot_3')
// (6, 4, 'neigh_op_tnl_3')
// (6, 5, 'neigh_op_lft_3')
// (6, 6, 'neigh_op_bnl_3')

reg n151 = 0;
// (4, 4, 'neigh_op_tnr_5')
// (4, 5, 'neigh_op_rgt_5')
// (4, 6, 'neigh_op_bnr_5')
// (5, 4, 'neigh_op_top_5')
// (5, 5, 'local_g1_5')
// (5, 5, 'lutff_0/in_0')
// (5, 5, 'lutff_5/out')
// (5, 6, 'neigh_op_bot_5')
// (6, 4, 'neigh_op_tnl_5')
// (6, 5, 'neigh_op_lft_5')
// (6, 6, 'neigh_op_bnl_5')

reg n152 = 0;
// (4, 4, 'neigh_op_tnr_6')
// (4, 5, 'neigh_op_rgt_6')
// (4, 6, 'neigh_op_bnr_6')
// (5, 4, 'neigh_op_top_6')
// (5, 5, 'local_g1_6')
// (5, 5, 'lutff_3/in_0')
// (5, 5, 'lutff_6/out')
// (5, 6, 'neigh_op_bot_6')
// (6, 4, 'neigh_op_tnl_6')
// (6, 5, 'neigh_op_lft_6')
// (6, 6, 'neigh_op_bnl_6')

reg n153 = 0;
// (4, 4, 'neigh_op_tnr_7')
// (4, 5, 'neigh_op_rgt_7')
// (4, 6, 'neigh_op_bnr_7')
// (5, 3, 'sp4_r_v_b_39')
// (5, 4, 'local_g0_2')
// (5, 4, 'lutff_6/in_0')
// (5, 4, 'neigh_op_top_7')
// (5, 4, 'sp4_r_v_b_26')
// (5, 5, 'lutff_7/out')
// (5, 5, 'sp4_r_v_b_15')
// (5, 6, 'neigh_op_bot_7')
// (5, 6, 'sp4_r_v_b_2')
// (6, 2, 'sp4_v_t_39')
// (6, 3, 'sp4_v_b_39')
// (6, 4, 'neigh_op_tnl_7')
// (6, 4, 'sp4_v_b_26')
// (6, 5, 'neigh_op_lft_7')
// (6, 5, 'sp4_v_b_15')
// (6, 6, 'neigh_op_bnl_7')
// (6, 6, 'sp4_v_b_2')

reg n154 = 0;
// (4, 5, 'neigh_op_tnr_1')
// (4, 6, 'neigh_op_rgt_1')
// (4, 7, 'neigh_op_bnr_1')
// (5, 5, 'neigh_op_top_1')
// (5, 6, 'local_g0_1')
// (5, 6, 'local_g1_1')
// (5, 6, 'lutff_0/in_0')
// (5, 6, 'lutff_1/out')
// (5, 6, 'lutff_4/in_1')
// (5, 7, 'neigh_op_bot_1')
// (6, 5, 'neigh_op_tnl_1')
// (6, 6, 'neigh_op_lft_1')
// (6, 7, 'neigh_op_bnl_1')

reg n155 = 0;
// (4, 5, 'neigh_op_tnr_3')
// (4, 6, 'neigh_op_rgt_3')
// (4, 7, 'neigh_op_bnr_3')
// (5, 5, 'neigh_op_top_3')
// (5, 6, 'local_g1_3')
// (5, 6, 'lutff_3/out')
// (5, 6, 'lutff_7/in_1')
// (5, 7, 'neigh_op_bot_3')
// (6, 5, 'neigh_op_tnl_3')
// (6, 6, 'neigh_op_lft_3')
// (6, 7, 'neigh_op_bnl_3')

reg n156 = 0;
// (4, 5, 'neigh_op_tnr_5')
// (4, 6, 'neigh_op_rgt_5')
// (4, 7, 'neigh_op_bnr_5')
// (5, 5, 'neigh_op_top_5')
// (5, 6, 'local_g0_5')
// (5, 6, 'lutff_3/in_2')
// (5, 6, 'lutff_5/out')
// (5, 6, 'lutff_6/in_1')
// (5, 7, 'neigh_op_bot_5')
// (6, 5, 'neigh_op_tnl_5')
// (6, 6, 'neigh_op_lft_5')
// (6, 7, 'neigh_op_bnl_5')

reg n157 = 0;
// (4, 5, 'neigh_op_tnr_6')
// (4, 6, 'neigh_op_rgt_6')
// (4, 7, 'neigh_op_bnr_6')
// (5, 5, 'neigh_op_top_6')
// (5, 6, 'local_g0_6')
// (5, 6, 'local_g1_6')
// (5, 6, 'lutff_1/in_1')
// (5, 6, 'lutff_6/out')
// (5, 6, 'lutff_7/in_2')
// (5, 7, 'neigh_op_bot_6')
// (6, 5, 'neigh_op_tnl_6')
// (6, 6, 'neigh_op_lft_6')
// (6, 7, 'neigh_op_bnl_6')

reg n158 = 0;
// (4, 5, 'neigh_op_tnr_7')
// (4, 6, 'neigh_op_rgt_7')
// (4, 7, 'neigh_op_bnr_7')
// (5, 5, 'neigh_op_top_7')
// (5, 6, 'local_g0_7')
// (5, 6, 'lutff_0/in_1')
// (5, 6, 'lutff_7/out')
// (5, 7, 'neigh_op_bot_7')
// (6, 5, 'neigh_op_tnl_7')
// (6, 6, 'neigh_op_lft_7')
// (6, 7, 'neigh_op_bnl_7')

wire n159;
// (4, 5, 'sp4_r_v_b_39')
// (4, 6, 'sp4_r_v_b_26')
// (4, 7, 'sp4_r_v_b_15')
// (4, 8, 'sp4_r_v_b_2')
// (5, 4, 'sp4_h_r_8')
// (5, 4, 'sp4_v_t_39')
// (5, 5, 'sp4_v_b_39')
// (5, 6, 'sp4_v_b_26')
// (5, 7, 'sp4_v_b_15')
// (5, 8, 'sp4_h_r_2')
// (5, 8, 'sp4_v_b_2')
// (6, 3, 'neigh_op_tnr_0')
// (6, 4, 'neigh_op_rgt_0')
// (6, 4, 'sp4_h_r_21')
// (6, 5, 'neigh_op_bnr_0')
// (6, 7, 'sp4_r_v_b_39')
// (6, 8, 'sp4_h_r_15')
// (6, 8, 'sp4_r_v_b_26')
// (6, 9, 'sp4_r_v_b_15')
// (6, 10, 'sp4_r_v_b_2')
// (7, 0, 'span12_vert_23')
// (7, 1, 'sp12_v_b_23')
// (7, 2, 'sp12_v_b_20')
// (7, 2, 'sp4_r_v_b_41')
// (7, 3, 'neigh_op_top_0')
// (7, 3, 'sp12_v_b_19')
// (7, 3, 'sp4_r_v_b_28')
// (7, 4, 'lutff_0/out')
// (7, 4, 'sp12_v_b_16')
// (7, 4, 'sp4_h_r_32')
// (7, 4, 'sp4_r_v_b_17')
// (7, 5, 'neigh_op_bot_0')
// (7, 5, 'sp12_v_b_15')
// (7, 5, 'sp4_r_v_b_4')
// (7, 6, 'sp12_v_b_12')
// (7, 6, 'sp4_r_v_b_41')
// (7, 6, 'sp4_v_t_39')
// (7, 7, 'sp12_v_b_11')
// (7, 7, 'sp4_r_v_b_28')
// (7, 7, 'sp4_v_b_39')
// (7, 8, 'sp12_v_b_8')
// (7, 8, 'sp4_h_r_26')
// (7, 8, 'sp4_r_v_b_17')
// (7, 8, 'sp4_v_b_26')
// (7, 9, 'local_g2_7')
// (7, 9, 'local_g3_7')
// (7, 9, 'lutff_5/in_1')
// (7, 9, 'lutff_6/in_1')
// (7, 9, 'sp12_v_b_7')
// (7, 9, 'sp4_r_v_b_4')
// (7, 9, 'sp4_v_b_15')
// (7, 10, 'local_g0_2')
// (7, 10, 'local_g1_2')
// (7, 10, 'lutff_2/in_3')
// (7, 10, 'lutff_3/in_1')
// (7, 10, 'sp12_v_b_4')
// (7, 10, 'sp4_h_r_8')
// (7, 10, 'sp4_r_v_b_37')
// (7, 10, 'sp4_v_b_2')
// (7, 11, 'sp12_v_b_3')
// (7, 11, 'sp4_r_v_b_24')
// (7, 12, 'sp12_v_b_0')
// (7, 12, 'sp4_r_v_b_13')
// (7, 13, 'sp4_r_v_b_0')
// (8, 1, 'sp4_v_t_41')
// (8, 2, 'sp4_v_b_41')
// (8, 3, 'neigh_op_tnl_0')
// (8, 3, 'sp4_v_b_28')
// (8, 4, 'neigh_op_lft_0')
// (8, 4, 'sp4_h_r_45')
// (8, 4, 'sp4_v_b_17')
// (8, 5, 'neigh_op_bnl_0')
// (8, 5, 'sp4_r_v_b_36')
// (8, 5, 'sp4_v_b_4')
// (8, 5, 'sp4_v_t_41')
// (8, 6, 'sp4_r_v_b_25')
// (8, 6, 'sp4_v_b_41')
// (8, 7, 'sp4_r_v_b_12')
// (8, 7, 'sp4_v_b_28')
// (8, 8, 'sp4_h_r_39')
// (8, 8, 'sp4_r_v_b_1')
// (8, 8, 'sp4_v_b_17')
// (8, 9, 'local_g0_4')
// (8, 9, 'lutff_0/in_0')
// (8, 9, 'lutff_1/in_1')
// (8, 9, 'sp4_r_v_b_36')
// (8, 9, 'sp4_r_v_b_39')
// (8, 9, 'sp4_v_b_4')
// (8, 9, 'sp4_v_t_37')
// (8, 10, 'sp4_h_r_21')
// (8, 10, 'sp4_r_v_b_25')
// (8, 10, 'sp4_r_v_b_26')
// (8, 10, 'sp4_v_b_37')
// (8, 11, 'local_g2_0')
// (8, 11, 'lutff_3/in_3')
// (8, 11, 'sp4_r_v_b_12')
// (8, 11, 'sp4_r_v_b_15')
// (8, 11, 'sp4_v_b_24')
// (8, 12, 'sp4_r_v_b_1')
// (8, 12, 'sp4_r_v_b_2')
// (8, 12, 'sp4_v_b_13')
// (8, 13, 'sp4_v_b_0')
// (9, 4, 'sp4_h_l_45')
// (9, 4, 'sp4_v_t_36')
// (9, 5, 'sp4_v_b_36')
// (9, 6, 'sp4_v_b_25')
// (9, 7, 'local_g0_4')
// (9, 7, 'lutff_0/in_2')
// (9, 7, 'sp4_v_b_12')
// (9, 8, 'sp4_h_l_39')
// (9, 8, 'sp4_v_b_1')
// (9, 8, 'sp4_v_t_36')
// (9, 8, 'sp4_v_t_39')
// (9, 9, 'sp4_v_b_36')
// (9, 9, 'sp4_v_b_39')
// (9, 10, 'local_g2_0')
// (9, 10, 'local_g3_0')
// (9, 10, 'lutff_1/in_3')
// (9, 10, 'lutff_7/in_2')
// (9, 10, 'sp4_h_r_32')
// (9, 10, 'sp4_v_b_25')
// (9, 10, 'sp4_v_b_26')
// (9, 11, 'local_g0_4')
// (9, 11, 'local_g0_7')
// (9, 11, 'lutff_2/in_3')
// (9, 11, 'lutff_6/in_2')
// (9, 11, 'sp4_v_b_12')
// (9, 11, 'sp4_v_b_15')
// (9, 12, 'sp4_v_b_1')
// (9, 12, 'sp4_v_b_2')
// (10, 10, 'sp4_h_r_45')
// (11, 10, 'sp4_h_l_45')

reg n160 = 0;
// (4, 5, 'sp4_r_v_b_40')
// (4, 6, 'local_g1_5')
// (4, 6, 'lutff_1/in_3')
// (4, 6, 'sp4_r_v_b_29')
// (4, 7, 'sp4_r_v_b_16')
// (4, 8, 'sp4_r_v_b_5')
// (5, 3, 'neigh_op_tnr_3')
// (5, 4, 'local_g3_3')
// (5, 4, 'lutff_2/in_2')
// (5, 4, 'neigh_op_rgt_3')
// (5, 4, 'sp4_h_r_11')
// (5, 4, 'sp4_v_t_40')
// (5, 5, 'neigh_op_bnr_3')
// (5, 5, 'sp4_v_b_40')
// (5, 6, 'sp4_v_b_29')
// (5, 7, 'sp4_v_b_16')
// (5, 8, 'sp4_v_b_5')
// (6, 3, 'neigh_op_top_3')
// (6, 4, 'local_g1_3')
// (6, 4, 'lutff_3/out')
// (6, 4, 'lutff_7/in_3')
// (6, 4, 'sp4_h_r_22')
// (6, 5, 'neigh_op_bot_3')
// (7, 3, 'neigh_op_tnl_3')
// (7, 4, 'neigh_op_lft_3')
// (7, 4, 'sp4_h_r_35')
// (7, 5, 'neigh_op_bnl_3')
// (8, 4, 'sp4_h_r_46')
// (9, 4, 'sp4_h_l_46')

reg n161 = 0;
// (4, 6, 'neigh_op_tnr_3')
// (4, 7, 'neigh_op_rgt_3')
// (4, 8, 'neigh_op_bnr_3')
// (5, 6, 'neigh_op_top_3')
// (5, 7, 'lutff_3/out')
// (5, 8, 'neigh_op_bot_3')
// (6, 6, 'neigh_op_tnl_3')
// (6, 7, 'local_g0_3')
// (6, 7, 'lutff_0/in_1')
// (6, 7, 'lutff_2/in_1')
// (6, 7, 'neigh_op_lft_3')
// (6, 8, 'neigh_op_bnl_3')

reg n162 = 0;
// (4, 6, 'neigh_op_tnr_4')
// (4, 7, 'neigh_op_rgt_4')
// (4, 8, 'neigh_op_bnr_4')
// (5, 6, 'neigh_op_top_4')
// (5, 7, 'local_g0_4')
// (5, 7, 'lutff_0/in_0')
// (5, 7, 'lutff_4/out')
// (5, 8, 'local_g1_4')
// (5, 8, 'lutff_7/in_0')
// (5, 8, 'neigh_op_bot_4')
// (6, 6, 'neigh_op_tnl_4')
// (6, 7, 'neigh_op_lft_4')
// (6, 8, 'neigh_op_bnl_4')

reg n163 = 0;
// (4, 6, 'neigh_op_tnr_5')
// (4, 7, 'neigh_op_rgt_5')
// (4, 7, 'sp4_r_v_b_42')
// (4, 8, 'neigh_op_bnr_5')
// (4, 8, 'sp4_r_v_b_31')
// (4, 9, 'sp4_r_v_b_18')
// (4, 10, 'sp4_r_v_b_7')
// (4, 11, 'sp4_r_v_b_42')
// (4, 12, 'sp4_r_v_b_31')
// (4, 13, 'sp4_r_v_b_18')
// (4, 14, 'sp4_r_v_b_7')
// (5, 6, 'neigh_op_top_5')
// (5, 6, 'sp4_v_t_42')
// (5, 7, 'lutff_5/out')
// (5, 7, 'sp4_v_b_42')
// (5, 8, 'neigh_op_bot_5')
// (5, 8, 'sp4_v_b_31')
// (5, 9, 'sp4_v_b_18')
// (5, 10, 'local_g1_7')
// (5, 10, 'lutff_4/in_0')
// (5, 10, 'sp4_v_b_7')
// (5, 10, 'sp4_v_t_42')
// (5, 11, 'local_g2_2')
// (5, 11, 'lutff_1/in_3')
// (5, 11, 'sp4_v_b_42')
// (5, 12, 'sp4_v_b_31')
// (5, 13, 'sp4_v_b_18')
// (5, 14, 'sp4_v_b_7')
// (6, 6, 'neigh_op_tnl_5')
// (6, 7, 'neigh_op_lft_5')
// (6, 8, 'neigh_op_bnl_5')

reg n164 = 0;
// (4, 6, 'neigh_op_tnr_6')
// (4, 7, 'neigh_op_rgt_6')
// (4, 8, 'neigh_op_bnr_6')
// (5, 6, 'neigh_op_top_6')
// (5, 7, 'local_g1_6')
// (5, 7, 'lutff_6/out')
// (5, 7, 'lutff_7/in_0')
// (5, 8, 'neigh_op_bot_6')
// (6, 6, 'neigh_op_tnl_6')
// (6, 7, 'neigh_op_lft_6')
// (6, 8, 'neigh_op_bnl_6')

reg n165 = 0;
// (4, 6, 'sp12_h_r_1')
// (5, 6, 'sp12_h_r_2')
// (6, 6, 'sp12_h_r_5')
// (7, 6, 'sp12_h_r_6')
// (8, 5, 'neigh_op_tnr_1')
// (8, 6, 'neigh_op_rgt_1')
// (8, 6, 'sp12_h_r_9')
// (8, 7, 'neigh_op_bnr_1')
// (9, 5, 'neigh_op_top_1')
// (9, 6, 'lutff_1/out')
// (9, 6, 'sp12_h_r_10')
// (9, 7, 'neigh_op_bot_1')
// (10, 5, 'neigh_op_tnl_1')
// (10, 6, 'neigh_op_lft_1')
// (10, 6, 'sp12_h_r_13')
// (10, 7, 'neigh_op_bnl_1')
// (11, 6, 'local_g0_6')
// (11, 6, 'lutff_6/in_0')
// (11, 6, 'sp12_h_r_14')
// (12, 6, 'sp12_h_r_17')
// (13, 6, 'span12_horz_17')

wire n166;
// (4, 6, 'sp4_r_v_b_37')
// (4, 7, 'sp4_r_v_b_24')
// (4, 8, 'neigh_op_tnr_0')
// (4, 8, 'sp4_r_v_b_13')
// (4, 9, 'neigh_op_rgt_0')
// (4, 9, 'sp4_r_v_b_0')
// (4, 10, 'neigh_op_bnr_0')
// (5, 5, 'sp4_v_t_37')
// (5, 6, 'local_g2_5')
// (5, 6, 'local_g3_5')
// (5, 6, 'lutff_4/in_3')
// (5, 6, 'lutff_5/in_3')
// (5, 6, 'sp4_v_b_37')
// (5, 7, 'sp4_v_b_24')
// (5, 8, 'neigh_op_top_0')
// (5, 8, 'sp4_v_b_13')
// (5, 9, 'local_g2_0')
// (5, 9, 'lutff_0/out')
// (5, 9, 'lutff_7/in_3')
// (5, 9, 'sp4_v_b_0')
// (5, 10, 'neigh_op_bot_0')
// (6, 8, 'neigh_op_tnl_0')
// (6, 9, 'neigh_op_lft_0')
// (6, 10, 'neigh_op_bnl_0')

wire n167;
// (4, 6, 'sp4_r_v_b_45')
// (4, 7, 'sp4_r_v_b_32')
// (4, 8, 'sp4_r_v_b_21')
// (4, 9, 'sp4_r_v_b_8')
// (5, 5, 'sp4_v_t_45')
// (5, 6, 'sp4_v_b_45')
// (5, 7, 'sp4_v_b_32')
// (5, 8, 'local_g0_5')
// (5, 8, 'lutff_7/in_2')
// (5, 8, 'sp4_v_b_21')
// (5, 9, 'sp4_h_r_8')
// (5, 9, 'sp4_v_b_8')
// (6, 3, 'sp4_r_v_b_36')
// (6, 4, 'local_g0_1')
// (6, 4, 'lutff_7/in_2')
// (6, 4, 'sp4_r_v_b_25')
// (6, 5, 'sp4_r_v_b_12')
// (6, 6, 'sp4_r_v_b_1')
// (6, 7, 'sp4_r_v_b_40')
// (6, 8, 'neigh_op_tnr_0')
// (6, 8, 'sp4_r_v_b_29')
// (6, 9, 'neigh_op_rgt_0')
// (6, 9, 'sp4_h_r_21')
// (6, 9, 'sp4_r_v_b_16')
// (6, 10, 'neigh_op_bnr_0')
// (6, 10, 'sp4_r_v_b_5')
// (7, 2, 'sp4_v_t_36')
// (7, 3, 'sp4_v_b_36')
// (7, 4, 'sp4_v_b_25')
// (7, 5, 'sp4_v_b_12')
// (7, 6, 'sp4_r_v_b_36')
// (7, 6, 'sp4_v_b_1')
// (7, 6, 'sp4_v_t_40')
// (7, 7, 'sp4_r_v_b_25')
// (7, 7, 'sp4_v_b_40')
// (7, 8, 'neigh_op_top_0')
// (7, 8, 'sp4_r_v_b_12')
// (7, 8, 'sp4_v_b_29')
// (7, 9, 'lutff_0/out')
// (7, 9, 'sp4_h_r_32')
// (7, 9, 'sp4_r_v_b_1')
// (7, 9, 'sp4_v_b_16')
// (7, 10, 'neigh_op_bot_0')
// (7, 10, 'sp4_v_b_5')
// (8, 5, 'sp4_v_t_36')
// (8, 6, 'sp4_v_b_36')
// (8, 7, 'local_g2_1')
// (8, 7, 'local_g3_1')
// (8, 7, 'lutff_2/in_3')
// (8, 7, 'lutff_3/in_2')
// (8, 7, 'lutff_7/in_3')
// (8, 7, 'sp4_v_b_25')
// (8, 8, 'neigh_op_tnl_0')
// (8, 8, 'sp4_v_b_12')
// (8, 9, 'neigh_op_lft_0')
// (8, 9, 'sp4_h_r_45')
// (8, 9, 'sp4_v_b_1')
// (8, 10, 'neigh_op_bnl_0')
// (9, 9, 'sp4_h_l_45')

wire n168;
// (4, 6, 'sp4_r_v_b_47')
// (4, 7, 'sp4_r_v_b_34')
// (4, 8, 'sp4_r_v_b_23')
// (4, 9, 'sp4_r_v_b_10')
// (5, 5, 'sp4_v_t_47')
// (5, 6, 'sp4_v_b_47')
// (5, 7, 'sp4_v_b_34')
// (5, 8, 'local_g0_7')
// (5, 8, 'lutff_5/in_2')
// (5, 8, 'sp4_v_b_23')
// (5, 9, 'sp4_h_r_10')
// (5, 9, 'sp4_v_b_10')
// (6, 8, 'neigh_op_tnr_1')
// (6, 9, 'neigh_op_rgt_1')
// (6, 9, 'sp4_h_r_23')
// (6, 10, 'neigh_op_bnr_1')
// (7, 8, 'neigh_op_top_1')
// (7, 9, 'local_g2_1')
// (7, 9, 'lutff_0/in_1')
// (7, 9, 'lutff_1/out')
// (7, 9, 'sp4_h_r_34')
// (7, 10, 'neigh_op_bot_1')
// (8, 8, 'neigh_op_tnl_1')
// (8, 9, 'neigh_op_lft_1')
// (8, 9, 'sp4_h_r_47')
// (8, 10, 'neigh_op_bnl_1')
// (9, 9, 'sp4_h_l_47')

reg n169 = 0;
// (4, 7, 'local_g3_1')
// (4, 7, 'lutff_6/in_0')
// (4, 7, 'sp4_r_v_b_41')
// (4, 8, 'sp4_r_v_b_28')
// (4, 8, 'sp4_r_v_b_44')
// (4, 9, 'neigh_op_tnr_2')
// (4, 9, 'sp4_r_v_b_17')
// (4, 9, 'sp4_r_v_b_33')
// (4, 10, 'local_g3_2')
// (4, 10, 'lutff_3/in_0')
// (4, 10, 'neigh_op_rgt_2')
// (4, 10, 'sp4_r_v_b_20')
// (4, 10, 'sp4_r_v_b_4')
// (4, 11, 'neigh_op_bnr_2')
// (4, 11, 'sp4_r_v_b_9')
// (5, 6, 'sp4_v_t_41')
// (5, 7, 'sp4_h_r_2')
// (5, 7, 'sp4_v_b_41')
// (5, 7, 'sp4_v_t_44')
// (5, 8, 'sp4_v_b_28')
// (5, 8, 'sp4_v_b_44')
// (5, 9, 'neigh_op_top_2')
// (5, 9, 'sp4_v_b_17')
// (5, 9, 'sp4_v_b_33')
// (5, 10, 'lutff_2/out')
// (5, 10, 'sp4_v_b_20')
// (5, 10, 'sp4_v_b_4')
// (5, 11, 'neigh_op_bot_2')
// (5, 11, 'sp4_v_b_9')
// (6, 7, 'sp4_h_r_15')
// (6, 9, 'neigh_op_tnl_2')
// (6, 10, 'neigh_op_lft_2')
// (6, 11, 'neigh_op_bnl_2')
// (7, 7, 'sp4_h_r_26')
// (8, 7, 'local_g2_7')
// (8, 7, 'lutff_0/in_3')
// (8, 7, 'sp4_h_r_39')
// (9, 7, 'sp4_h_l_39')

reg n170 = 0;
// (4, 7, 'neigh_op_tnr_0')
// (4, 8, 'neigh_op_rgt_0')
// (4, 9, 'neigh_op_bnr_0')
// (5, 7, 'neigh_op_top_0')
// (5, 8, 'local_g0_0')
// (5, 8, 'lutff_0/out')
// (5, 8, 'lutff_4/in_0')
// (5, 9, 'neigh_op_bot_0')
// (6, 7, 'neigh_op_tnl_0')
// (6, 8, 'neigh_op_lft_0')
// (6, 9, 'neigh_op_bnl_0')

reg n171 = 0;
// (4, 7, 'neigh_op_tnr_1')
// (4, 8, 'neigh_op_rgt_1')
// (4, 9, 'neigh_op_bnr_1')
// (5, 7, 'neigh_op_top_1')
// (5, 8, 'local_g1_1')
// (5, 8, 'lutff_1/out')
// (5, 8, 'lutff_6/in_0')
// (5, 9, 'neigh_op_bot_1')
// (6, 7, 'neigh_op_tnl_1')
// (6, 8, 'neigh_op_lft_1')
// (6, 9, 'neigh_op_bnl_1')

reg n172 = 0;
// (4, 7, 'neigh_op_tnr_2')
// (4, 8, 'neigh_op_rgt_2')
// (4, 9, 'neigh_op_bnr_2')
// (5, 7, 'neigh_op_top_2')
// (5, 8, 'local_g1_2')
// (5, 8, 'lutff_2/out')
// (5, 8, 'lutff_3/in_0')
// (5, 9, 'neigh_op_bot_2')
// (6, 7, 'neigh_op_tnl_2')
// (6, 8, 'neigh_op_lft_2')
// (6, 9, 'neigh_op_bnl_2')

reg n173 = 0;
// (4, 7, 'neigh_op_tnr_3')
// (4, 8, 'neigh_op_rgt_3')
// (4, 8, 'sp4_r_v_b_38')
// (4, 9, 'neigh_op_bnr_3')
// (4, 9, 'sp4_r_v_b_27')
// (4, 10, 'sp4_r_v_b_14')
// (4, 11, 'sp4_r_v_b_3')
// (5, 7, 'neigh_op_top_3')
// (5, 7, 'sp4_v_t_38')
// (5, 8, 'lutff_3/out')
// (5, 8, 'sp4_v_b_38')
// (5, 9, 'neigh_op_bot_3')
// (5, 9, 'sp4_v_b_27')
// (5, 10, 'local_g1_6')
// (5, 10, 'lutff_6/in_3')
// (5, 10, 'sp4_v_b_14')
// (5, 11, 'sp4_v_b_3')
// (6, 7, 'neigh_op_tnl_3')
// (6, 8, 'neigh_op_lft_3')
// (6, 9, 'neigh_op_bnl_3')

reg n174 = 0;
// (4, 7, 'neigh_op_tnr_4')
// (4, 8, 'neigh_op_rgt_4')
// (4, 9, 'neigh_op_bnr_4')
// (5, 7, 'neigh_op_top_4')
// (5, 8, 'local_g3_4')
// (5, 8, 'lutff_1/in_0')
// (5, 8, 'lutff_4/out')
// (5, 9, 'neigh_op_bot_4')
// (6, 7, 'neigh_op_tnl_4')
// (6, 8, 'neigh_op_lft_4')
// (6, 9, 'neigh_op_bnl_4')

reg n175 = 0;
// (4, 7, 'neigh_op_tnr_6')
// (4, 8, 'neigh_op_rgt_6')
// (4, 9, 'neigh_op_bnr_6')
// (5, 7, 'neigh_op_top_6')
// (5, 8, 'local_g0_6')
// (5, 8, 'lutff_2/in_0')
// (5, 8, 'lutff_6/out')
// (5, 9, 'neigh_op_bot_6')
// (6, 7, 'neigh_op_tnl_6')
// (6, 8, 'neigh_op_lft_6')
// (6, 9, 'neigh_op_bnl_6')

reg n176 = 0;
// (4, 7, 'sp4_r_v_b_45')
// (4, 8, 'sp4_r_v_b_32')
// (4, 9, 'neigh_op_tnr_4')
// (4, 9, 'sp4_r_v_b_21')
// (4, 10, 'local_g2_4')
// (4, 10, 'lutff_6/in_0')
// (4, 10, 'neigh_op_rgt_4')
// (4, 10, 'sp4_r_v_b_8')
// (4, 11, 'neigh_op_bnr_4')
// (5, 6, 'sp4_v_t_45')
// (5, 7, 'sp4_r_v_b_44')
// (5, 7, 'sp4_v_b_45')
// (5, 8, 'sp4_r_v_b_33')
// (5, 8, 'sp4_v_b_32')
// (5, 9, 'local_g1_5')
// (5, 9, 'lutff_1/in_3')
// (5, 9, 'neigh_op_top_4')
// (5, 9, 'sp4_r_v_b_20')
// (5, 9, 'sp4_v_b_21')
// (5, 10, 'lutff_4/out')
// (5, 10, 'sp4_r_v_b_9')
// (5, 10, 'sp4_v_b_8')
// (5, 11, 'neigh_op_bot_4')
// (6, 6, 'sp4_v_t_44')
// (6, 7, 'sp4_v_b_44')
// (6, 8, 'local_g3_1')
// (6, 8, 'lutff_0/in_0')
// (6, 8, 'sp4_v_b_33')
// (6, 9, 'neigh_op_tnl_4')
// (6, 9, 'sp4_v_b_20')
// (6, 10, 'neigh_op_lft_4')
// (6, 10, 'sp4_v_b_9')
// (6, 11, 'neigh_op_bnl_4')

reg n177 = 0;
// (4, 8, 'neigh_op_tnr_2')
// (4, 9, 'neigh_op_rgt_2')
// (4, 10, 'neigh_op_bnr_2')
// (5, 8, 'neigh_op_top_2')
// (5, 9, 'local_g0_2')
// (5, 9, 'local_g1_2')
// (5, 9, 'lutff_1/in_0')
// (5, 9, 'lutff_2/out')
// (5, 9, 'lutff_3/in_1')
// (5, 10, 'neigh_op_bot_2')
// (6, 8, 'neigh_op_tnl_2')
// (6, 9, 'neigh_op_lft_2')
// (6, 10, 'neigh_op_bnl_2')

reg n178 = 0;
// (4, 8, 'neigh_op_tnr_3')
// (4, 9, 'local_g2_3')
// (4, 9, 'lutff_7/in_0')
// (4, 9, 'neigh_op_rgt_3')
// (4, 10, 'neigh_op_bnr_3')
// (5, 8, 'neigh_op_top_3')
// (5, 9, 'local_g2_3')
// (5, 9, 'lutff_3/out')
// (5, 9, 'lutff_7/in_2')
// (5, 10, 'neigh_op_bot_3')
// (6, 8, 'neigh_op_tnl_3')
// (6, 9, 'neigh_op_lft_3')
// (6, 10, 'neigh_op_bnl_3')

reg n179 = 0;
// (4, 8, 'neigh_op_tnr_4')
// (4, 9, 'neigh_op_rgt_4')
// (4, 10, 'neigh_op_bnr_4')
// (5, 8, 'neigh_op_top_4')
// (5, 9, 'local_g2_4')
// (5, 9, 'local_g3_4')
// (5, 9, 'lutff_2/in_1')
// (5, 9, 'lutff_4/out')
// (5, 9, 'lutff_6/in_2')
// (5, 10, 'neigh_op_bot_4')
// (6, 8, 'neigh_op_tnl_4')
// (6, 9, 'neigh_op_lft_4')
// (6, 10, 'neigh_op_bnl_4')

reg n180 = 0;
// (4, 8, 'neigh_op_tnr_5')
// (4, 9, 'neigh_op_rgt_5')
// (4, 10, 'neigh_op_bnr_5')
// (5, 8, 'neigh_op_top_5')
// (5, 9, 'local_g0_5')
// (5, 9, 'lutff_5/out')
// (5, 9, 'lutff_6/in_1')
// (5, 10, 'neigh_op_bot_5')
// (6, 8, 'neigh_op_tnl_5')
// (6, 9, 'neigh_op_lft_5')
// (6, 10, 'neigh_op_bnl_5')

reg n181 = 0;
// (4, 8, 'neigh_op_tnr_6')
// (4, 9, 'neigh_op_rgt_6')
// (4, 10, 'neigh_op_bnr_6')
// (5, 8, 'neigh_op_top_6')
// (5, 9, 'local_g0_6')
// (5, 9, 'lutff_1/in_1')
// (5, 9, 'lutff_6/out')
// (5, 10, 'neigh_op_bot_6')
// (6, 8, 'neigh_op_tnl_6')
// (6, 9, 'neigh_op_lft_6')
// (6, 10, 'neigh_op_bnl_6')

reg n182 = 0;
// (4, 8, 'neigh_op_tnr_7')
// (4, 9, 'neigh_op_rgt_7')
// (4, 10, 'neigh_op_bnr_7')
// (5, 8, 'neigh_op_top_7')
// (5, 9, 'local_g0_7')
// (5, 9, 'lutff_4/in_1')
// (5, 9, 'lutff_5/in_2')
// (5, 9, 'lutff_7/out')
// (5, 10, 'neigh_op_bot_7')
// (6, 8, 'neigh_op_tnl_7')
// (6, 9, 'neigh_op_lft_7')
// (6, 10, 'neigh_op_bnl_7')

reg n183 = 0;
// (4, 8, 'sp4_r_v_b_36')
// (4, 9, 'neigh_op_tnr_6')
// (4, 9, 'sp4_r_v_b_25')
// (4, 10, 'neigh_op_rgt_6')
// (4, 10, 'sp4_r_v_b_12')
// (4, 11, 'local_g1_1')
// (4, 11, 'lutff_6/in_0')
// (4, 11, 'neigh_op_bnr_6')
// (4, 11, 'sp4_r_v_b_1')
// (5, 7, 'sp4_v_t_36')
// (5, 8, 'sp4_v_b_36')
// (5, 9, 'neigh_op_top_6')
// (5, 9, 'sp4_v_b_25')
// (5, 10, 'lutff_6/out')
// (5, 10, 'sp4_v_b_12')
// (5, 11, 'neigh_op_bot_6')
// (5, 11, 'sp4_v_b_1')
// (6, 9, 'neigh_op_tnl_6')
// (6, 10, 'neigh_op_lft_6')
// (6, 11, 'neigh_op_bnl_6')

reg n184 = 0;
// (4, 9, 'neigh_op_tnr_0')
// (4, 9, 'sp4_r_v_b_45')
// (4, 10, 'neigh_op_rgt_0')
// (4, 10, 'sp4_r_v_b_32')
// (4, 11, 'neigh_op_bnr_0')
// (4, 11, 'sp4_r_v_b_21')
// (4, 12, 'sp4_r_v_b_8')
// (5, 0, 'span12_vert_19')
// (5, 1, 'sp12_v_b_19')
// (5, 2, 'sp12_v_b_16')
// (5, 3, 'local_g2_7')
// (5, 3, 'lutff_5/in_0')
// (5, 3, 'sp12_v_b_15')
// (5, 3, 'sp4_r_v_b_41')
// (5, 4, 'sp12_v_b_12')
// (5, 4, 'sp4_r_v_b_28')
// (5, 5, 'sp12_v_b_11')
// (5, 5, 'sp4_r_v_b_17')
// (5, 6, 'sp12_v_b_8')
// (5, 6, 'sp4_r_v_b_4')
// (5, 7, 'sp12_v_b_7')
// (5, 7, 'sp4_r_v_b_36')
// (5, 8, 'sp12_v_b_4')
// (5, 8, 'sp4_r_v_b_25')
// (5, 8, 'sp4_v_t_45')
// (5, 9, 'neigh_op_top_0')
// (5, 9, 'sp12_v_b_3')
// (5, 9, 'sp4_r_v_b_12')
// (5, 9, 'sp4_v_b_45')
// (5, 10, 'lutff_0/out')
// (5, 10, 'sp12_v_b_0')
// (5, 10, 'sp4_r_v_b_1')
// (5, 10, 'sp4_v_b_32')
// (5, 11, 'neigh_op_bot_0')
// (5, 11, 'sp4_v_b_21')
// (5, 12, 'local_g0_0')
// (5, 12, 'lutff_6/in_0')
// (5, 12, 'sp4_v_b_8')
// (6, 2, 'sp4_v_t_41')
// (6, 3, 'local_g2_1')
// (6, 3, 'lutff_0/in_3')
// (6, 3, 'sp4_v_b_41')
// (6, 4, 'sp4_v_b_28')
// (6, 5, 'sp4_v_b_17')
// (6, 6, 'sp4_v_b_4')
// (6, 6, 'sp4_v_t_36')
// (6, 7, 'sp4_v_b_36')
// (6, 8, 'sp4_v_b_25')
// (6, 9, 'neigh_op_tnl_0')
// (6, 9, 'sp4_v_b_12')
// (6, 10, 'neigh_op_lft_0')
// (6, 10, 'sp4_v_b_1')
// (6, 11, 'neigh_op_bnl_0')

reg n185 = 0;
// (4, 9, 'neigh_op_tnr_1')
// (4, 10, 'neigh_op_rgt_1')
// (4, 11, 'neigh_op_bnr_1')
// (5, 0, 'span12_vert_21')
// (5, 1, 'sp12_v_b_21')
// (5, 2, 'sp12_v_b_18')
// (5, 3, 'sp12_v_b_17')
// (5, 4, 'sp12_v_b_14')
// (5, 5, 'sp12_v_b_13')
// (5, 6, 'sp12_v_b_10')
// (5, 7, 'sp12_v_b_9')
// (5, 8, 'sp12_v_b_6')
// (5, 9, 'neigh_op_top_1')
// (5, 9, 'sp12_v_b_5')
// (5, 10, 'local_g1_1')
// (5, 10, 'lutff_0/in_0')
// (5, 10, 'lutff_1/out')
// (5, 10, 'sp12_v_b_2')
// (5, 11, 'local_g2_1')
// (5, 11, 'lutff_4/in_3')
// (5, 11, 'neigh_op_bot_1')
// (5, 11, 'sp12_v_b_1')
// (6, 9, 'neigh_op_tnl_1')
// (6, 10, 'neigh_op_lft_1')
// (6, 11, 'neigh_op_bnl_1')

reg \d_out[4] = 0 ;
// (4, 9, 'neigh_op_tnr_5')
// (4, 10, 'neigh_op_rgt_5')
// (4, 11, 'neigh_op_bnr_5')
// (5, 0, 'io_1/D_OUT_0')
// (5, 0, 'io_1/PAD')
// (5, 0, 'local_g0_5')
// (5, 0, 'span12_vert_5')
// (5, 1, 'sp12_v_b_5')
// (5, 2, 'sp12_v_b_2')
// (5, 3, 'sp12_v_b_1')
// (5, 3, 'sp12_v_t_22')
// (5, 4, 'sp12_v_b_22')
// (5, 5, 'sp12_v_b_21')
// (5, 6, 'sp12_v_b_18')
// (5, 7, 'sp12_v_b_17')
// (5, 8, 'sp12_v_b_14')
// (5, 9, 'neigh_op_top_5')
// (5, 9, 'sp12_v_b_13')
// (5, 10, 'lutff_5/out')
// (5, 10, 'sp12_v_b_10')
// (5, 11, 'neigh_op_bot_5')
// (5, 11, 'sp12_v_b_9')
// (5, 12, 'sp12_v_b_6')
// (5, 13, 'sp12_v_b_5')
// (5, 14, 'sp12_v_b_2')
// (5, 15, 'sp12_v_b_1')
// (6, 9, 'neigh_op_tnl_5')
// (6, 10, 'neigh_op_lft_5')
// (6, 11, 'neigh_op_bnl_5')

reg n187 = 0;
// (4, 9, 'sp12_h_r_1')
// (5, 9, 'sp12_h_r_2')
// (6, 9, 'sp12_h_r_5')
// (7, 9, 'sp12_h_r_6')
// (8, 9, 'sp12_h_r_9')
// (9, 9, 'local_g0_2')
// (9, 9, 'lutff_6/in_0')
// (9, 9, 'sp12_h_r_10')
// (10, 8, 'neigh_op_tnr_3')
// (10, 9, 'neigh_op_rgt_3')
// (10, 9, 'sp12_h_r_13')
// (10, 10, 'neigh_op_bnr_3')
// (11, 8, 'neigh_op_top_3')
// (11, 9, 'lutff_3/out')
// (11, 9, 'sp12_h_r_14')
// (11, 10, 'neigh_op_bot_3')
// (12, 8, 'neigh_op_tnl_3')
// (12, 9, 'neigh_op_lft_3')
// (12, 9, 'sp12_h_r_17')
// (12, 10, 'neigh_op_bnl_3')
// (13, 9, 'span12_horz_17')

reg n188 = 0;
// (4, 9, 'sp4_h_r_1')
// (5, 9, 'sp4_h_r_12')
// (6, 9, 'sp4_h_r_25')
// (7, 9, 'sp4_h_r_36')
// (7, 10, 'sp4_r_v_b_42')
// (7, 10, 'sp4_r_v_b_43')
// (7, 11, 'sp4_r_v_b_30')
// (7, 11, 'sp4_r_v_b_31')
// (7, 12, 'local_g1_1')
// (7, 12, 'lutff_5/in_1')
// (7, 12, 'lutff_7/in_1')
// (7, 12, 'sp4_h_r_1')
// (7, 12, 'sp4_r_v_b_18')
// (7, 12, 'sp4_r_v_b_19')
// (7, 13, 'sp4_r_v_b_6')
// (7, 13, 'sp4_r_v_b_7')
// (8, 9, 'sp4_h_l_36')
// (8, 9, 'sp4_v_t_42')
// (8, 9, 'sp4_v_t_43')
// (8, 10, 'sp4_v_b_42')
// (8, 10, 'sp4_v_b_43')
// (8, 11, 'sp4_v_b_30')
// (8, 11, 'sp4_v_b_31')
// (8, 12, 'local_g0_2')
// (8, 12, 'local_g1_4')
// (8, 12, 'lutff_1/in_1')
// (8, 12, 'lutff_2/in_2')
// (8, 12, 'lutff_5/in_2')
// (8, 12, 'lutff_6/in_1')
// (8, 12, 'sp4_h_r_12')
// (8, 12, 'sp4_v_b_18')
// (8, 12, 'sp4_v_b_19')
// (8, 13, 'local_g0_6')
// (8, 13, 'lutff_3/in_1')
// (8, 13, 'sp4_h_r_7')
// (8, 13, 'sp4_v_b_6')
// (8, 13, 'sp4_v_b_7')
// (9, 12, 'local_g2_1')
// (9, 12, 'lutff_1/in_2')
// (9, 12, 'sp4_h_r_25')
// (9, 13, 'local_g1_2')
// (9, 13, 'lutff_0/in_1')
// (9, 13, 'sp4_h_r_18')
// (10, 12, 'neigh_op_tnr_5')
// (10, 12, 'sp4_h_r_36')
// (10, 13, 'neigh_op_rgt_5')
// (10, 13, 'sp4_h_r_31')
// (10, 13, 'sp4_r_v_b_42')
// (10, 14, 'neigh_op_bnr_5')
// (10, 14, 'sp4_r_v_b_31')
// (10, 15, 'sp4_r_v_b_18')
// (10, 16, 'sp4_r_v_b_7')
// (11, 12, 'local_g0_5')
// (11, 12, 'lutff_1/in_0')
// (11, 12, 'neigh_op_top_5')
// (11, 12, 'sp4_h_l_36')
// (11, 12, 'sp4_v_t_42')
// (11, 13, 'local_g0_5')
// (11, 13, 'lutff_5/in_2')
// (11, 13, 'lutff_5/out')
// (11, 13, 'sp4_h_r_42')
// (11, 13, 'sp4_v_b_42')
// (11, 14, 'neigh_op_bot_5')
// (11, 14, 'sp4_v_b_31')
// (11, 15, 'sp4_v_b_18')
// (11, 16, 'sp4_v_b_7')
// (12, 12, 'neigh_op_tnl_5')
// (12, 13, 'neigh_op_lft_5')
// (12, 13, 'sp4_h_l_42')
// (12, 14, 'neigh_op_bnl_5')

wire n189;
// (4, 9, 'sp4_r_v_b_46')
// (4, 10, 'sp4_r_v_b_35')
// (4, 11, 'sp4_r_v_b_22')
// (4, 12, 'sp4_r_v_b_11')
// (4, 13, 'neigh_op_tnr_7')
// (4, 14, 'neigh_op_rgt_7')
// (4, 15, 'neigh_op_bnr_7')
// (5, 4, 'local_g3_7')
// (5, 4, 'lutff_0/in_0')
// (5, 4, 'lutff_2/in_0')
// (5, 4, 'lutff_3/in_1')
// (5, 4, 'sp4_r_v_b_47')
// (5, 5, 'sp4_r_v_b_34')
// (5, 6, 'sp4_r_v_b_23')
// (5, 7, 'sp4_r_v_b_10')
// (5, 8, 'sp4_h_r_11')
// (5, 8, 'sp4_h_r_4')
// (5, 8, 'sp4_r_v_b_39')
// (5, 8, 'sp4_v_t_46')
// (5, 9, 'sp12_v_t_22')
// (5, 9, 'sp4_r_v_b_26')
// (5, 9, 'sp4_v_b_46')
// (5, 10, 'local_g3_6')
// (5, 10, 'lutff_6/in_1')
// (5, 10, 'sp12_v_b_22')
// (5, 10, 'sp4_r_v_b_15')
// (5, 10, 'sp4_v_b_35')
// (5, 11, 'sp12_v_b_21')
// (5, 11, 'sp4_r_v_b_2')
// (5, 11, 'sp4_v_b_22')
// (5, 12, 'sp12_v_b_18')
// (5, 12, 'sp4_r_v_b_39')
// (5, 12, 'sp4_v_b_11')
// (5, 13, 'neigh_op_top_7')
// (5, 13, 'sp12_v_b_17')
// (5, 13, 'sp4_r_v_b_26')
// (5, 14, 'lutff_7/out')
// (5, 14, 'sp12_v_b_14')
// (5, 14, 'sp4_r_v_b_15')
// (5, 15, 'neigh_op_bot_7')
// (5, 15, 'sp12_v_b_13')
// (5, 15, 'sp4_r_v_b_2')
// (5, 16, 'sp12_v_b_10')
// (5, 17, 'span12_vert_9')
// (6, 3, 'sp4_v_t_47')
// (6, 4, 'sp4_v_b_47')
// (6, 5, 'sp4_v_b_34')
// (6, 6, 'sp4_v_b_23')
// (6, 7, 'sp4_v_b_10')
// (6, 7, 'sp4_v_t_39')
// (6, 8, 'sp4_h_r_17')
// (6, 8, 'sp4_h_r_22')
// (6, 8, 'sp4_v_b_39')
// (6, 9, 'sp4_v_b_26')
// (6, 10, 'local_g0_7')
// (6, 10, 'lutff_5/in_0')
// (6, 10, 'sp4_v_b_15')
// (6, 11, 'sp4_v_b_2')
// (6, 11, 'sp4_v_t_39')
// (6, 12, 'sp4_v_b_39')
// (6, 13, 'neigh_op_tnl_7')
// (6, 13, 'sp4_v_b_26')
// (6, 14, 'neigh_op_lft_7')
// (6, 14, 'sp4_v_b_15')
// (6, 15, 'local_g2_7')
// (6, 15, 'lutff_4/in_3')
// (6, 15, 'neigh_op_bnl_7')
// (6, 15, 'sp4_v_b_2')
// (7, 8, 'sp4_h_r_28')
// (7, 8, 'sp4_h_r_35')
// (8, 1, 'sp4_r_v_b_47')
// (8, 2, 'sp4_r_v_b_34')
// (8, 3, 'sp4_r_v_b_23')
// (8, 4, 'sp4_r_v_b_10')
// (8, 5, 'sp4_r_v_b_47')
// (8, 6, 'local_g0_1')
// (8, 6, 'lutff_6/in_1')
// (8, 6, 'sp4_r_v_b_34')
// (8, 7, 'sp4_r_v_b_23')
// (8, 8, 'local_g2_6')
// (8, 8, 'lutff_6/in_0')
// (8, 8, 'sp4_h_r_41')
// (8, 8, 'sp4_h_r_46')
// (8, 8, 'sp4_r_v_b_10')
// (9, 0, 'span4_vert_47')
// (9, 1, 'sp4_v_b_47')
// (9, 2, 'sp4_v_b_34')
// (9, 3, 'sp4_v_b_23')
// (9, 4, 'local_g0_2')
// (9, 4, 'lutff_0/in_0')
// (9, 4, 'sp4_v_b_10')
// (9, 4, 'sp4_v_t_47')
// (9, 5, 'sp4_v_b_47')
// (9, 6, 'sp4_v_b_34')
// (9, 7, 'sp4_v_b_23')
// (9, 8, 'sp4_h_l_41')
// (9, 8, 'sp4_h_l_46')
// (9, 8, 'sp4_v_b_10')

wire n190;
// (4, 10, 'neigh_op_tnr_0')
// (4, 11, 'neigh_op_rgt_0')
// (4, 12, 'neigh_op_bnr_0')
// (5, 10, 'neigh_op_top_0')
// (5, 11, 'lutff_0/out')
// (5, 12, 'neigh_op_bot_0')
// (6, 10, 'neigh_op_tnl_0')
// (6, 11, 'neigh_op_lft_0')
// (6, 12, 'local_g2_0')
// (6, 12, 'lutff_0/in_2')
// (6, 12, 'lutff_2/in_2')
// (6, 12, 'neigh_op_bnl_0')

wire n191;
// (4, 10, 'neigh_op_tnr_1')
// (4, 11, 'neigh_op_rgt_1')
// (4, 12, 'neigh_op_bnr_1')
// (5, 10, 'neigh_op_top_1')
// (5, 11, 'lutff_1/out')
// (5, 12, 'local_g0_1')
// (5, 12, 'lutff_3/in_0')
// (5, 12, 'neigh_op_bot_1')
// (6, 10, 'neigh_op_tnl_1')
// (6, 11, 'local_g1_1')
// (6, 11, 'lutff_2/in_0')
// (6, 11, 'neigh_op_lft_1')
// (6, 12, 'local_g2_1')
// (6, 12, 'lutff_7/in_2')
// (6, 12, 'neigh_op_bnl_1')

wire n192;
// (4, 10, 'neigh_op_tnr_3')
// (4, 11, 'neigh_op_rgt_3')
// (4, 12, 'neigh_op_bnr_3')
// (5, 10, 'neigh_op_top_3')
// (5, 11, 'lutff_3/out')
// (5, 12, 'local_g1_3')
// (5, 12, 'lutff_3/in_3')
// (5, 12, 'neigh_op_bot_3')
// (6, 10, 'neigh_op_tnl_3')
// (6, 11, 'local_g0_3')
// (6, 11, 'lutff_2/in_3')
// (6, 11, 'neigh_op_lft_3')
// (6, 12, 'local_g3_3')
// (6, 12, 'lutff_7/in_3')
// (6, 12, 'neigh_op_bnl_3')

wire n193;
// (4, 10, 'neigh_op_tnr_4')
// (4, 11, 'neigh_op_rgt_4')
// (4, 12, 'neigh_op_bnr_4')
// (5, 10, 'neigh_op_top_4')
// (5, 11, 'lutff_4/out')
// (5, 12, 'local_g0_4')
// (5, 12, 'lutff_3/in_1')
// (5, 12, 'lutff_4/in_2')
// (5, 12, 'neigh_op_bot_4')
// (6, 10, 'neigh_op_tnl_4')
// (6, 11, 'neigh_op_lft_4')
// (6, 12, 'neigh_op_bnl_4')

reg n194 = 0;
// (4, 10, 'neigh_op_tnr_6')
// (4, 11, 'local_g3_6')
// (4, 11, 'lutff_5/in_0')
// (4, 11, 'neigh_op_rgt_6')
// (4, 12, 'neigh_op_bnr_6')
// (5, 10, 'neigh_op_top_6')
// (5, 11, 'lutff_6/out')
// (5, 12, 'neigh_op_bot_6')
// (6, 10, 'neigh_op_tnl_6')
// (6, 11, 'neigh_op_lft_6')
// (6, 12, 'neigh_op_bnl_6')

wire n195;
// (4, 10, 'sp4_r_v_b_46')
// (4, 11, 'sp4_r_v_b_35')
// (4, 12, 'sp4_r_v_b_22')
// (4, 13, 'sp4_r_v_b_11')
// (5, 9, 'sp4_v_t_46')
// (5, 10, 'sp4_v_b_46')
// (5, 11, 'sp4_v_b_35')
// (5, 12, 'local_g0_6')
// (5, 12, 'lutff_5/in_1')
// (5, 12, 'sp4_v_b_22')
// (5, 13, 'sp4_h_r_6')
// (5, 13, 'sp4_v_b_11')
// (6, 12, 'neigh_op_tnr_7')
// (6, 13, 'neigh_op_rgt_7')
// (6, 13, 'sp4_h_r_19')
// (6, 14, 'neigh_op_bnr_7')
// (7, 12, 'local_g0_7')
// (7, 12, 'local_g1_7')
// (7, 12, 'lutff_2/in_0')
// (7, 12, 'lutff_3/in_0')
// (7, 12, 'lutff_6/in_1')
// (7, 12, 'neigh_op_top_7')
// (7, 13, 'lutff_7/out')
// (7, 13, 'sp4_h_r_30')
// (7, 14, 'neigh_op_bot_7')
// (8, 12, 'neigh_op_tnl_7')
// (8, 13, 'neigh_op_lft_7')
// (8, 13, 'sp4_h_r_43')
// (8, 14, 'neigh_op_bnl_7')
// (9, 13, 'sp4_h_l_43')

wire n196;
// (4, 11, 'neigh_op_tnr_0')
// (4, 12, 'neigh_op_rgt_0')
// (4, 13, 'neigh_op_bnr_0')
// (5, 11, 'neigh_op_top_0')
// (5, 12, 'local_g1_0')
// (5, 12, 'lutff_0/out')
// (5, 12, 'lutff_3/in_2')
// (5, 12, 'lutff_4/in_3')
// (5, 13, 'neigh_op_bot_0')
// (6, 11, 'neigh_op_tnl_0')
// (6, 12, 'neigh_op_lft_0')
// (6, 13, 'neigh_op_bnl_0')

wire n197;
// (4, 11, 'neigh_op_tnr_1')
// (4, 12, 'neigh_op_rgt_1')
// (4, 13, 'neigh_op_bnr_1')
// (5, 11, 'neigh_op_top_1')
// (5, 12, 'lutff_1/out')
// (5, 13, 'neigh_op_bot_1')
// (6, 11, 'neigh_op_tnl_1')
// (6, 12, 'local_g0_1')
// (6, 12, 'lutff_0/in_1')
// (6, 12, 'lutff_2/in_1')
// (6, 12, 'neigh_op_lft_1')
// (6, 13, 'neigh_op_bnl_1')

wire n198;
// (4, 11, 'neigh_op_tnr_3')
// (4, 12, 'neigh_op_rgt_3')
// (4, 13, 'neigh_op_bnr_3')
// (5, 11, 'neigh_op_top_3')
// (5, 12, 'lutff_3/out')
// (5, 13, 'neigh_op_bot_3')
// (6, 11, 'neigh_op_tnl_3')
// (6, 12, 'neigh_op_lft_3')
// (6, 13, 'local_g3_3')
// (6, 13, 'lutff_0/in_2')
// (6, 13, 'lutff_2/in_2')
// (6, 13, 'lutff_5/in_1')
// (6, 13, 'lutff_7/in_1')
// (6, 13, 'neigh_op_bnl_3')

wire n199;
// (4, 11, 'neigh_op_tnr_4')
// (4, 12, 'neigh_op_rgt_4')
// (4, 13, 'neigh_op_bnr_4')
// (5, 11, 'neigh_op_top_4')
// (5, 12, 'lutff_4/out')
// (5, 13, 'neigh_op_bot_4')
// (6, 11, 'neigh_op_tnl_4')
// (6, 12, 'local_g0_4')
// (6, 12, 'local_g1_4')
// (6, 12, 'lutff_4/in_1')
// (6, 12, 'lutff_5/in_1')
// (6, 12, 'lutff_6/in_0')
// (6, 12, 'neigh_op_lft_4')
// (6, 13, 'neigh_op_bnl_4')

reg n200 = 0;
// (4, 11, 'neigh_op_tnr_6')
// (4, 12, 'neigh_op_rgt_6')
// (4, 13, 'neigh_op_bnr_6')
// (5, 11, 'neigh_op_top_6')
// (5, 12, 'local_g1_6')
// (5, 12, 'lutff_0/in_3')
// (5, 12, 'lutff_6/out')
// (5, 13, 'neigh_op_bot_6')
// (6, 11, 'neigh_op_tnl_6')
// (6, 12, 'neigh_op_lft_6')
// (6, 13, 'neigh_op_bnl_6')

wire n201;
// (4, 11, 'sp12_h_r_1')
// (5, 11, 'sp12_h_r_2')
// (6, 11, 'sp12_h_r_5')
// (7, 11, 'local_g0_6')
// (7, 11, 'local_g1_6')
// (7, 11, 'lutff_0/in_0')
// (7, 11, 'lutff_1/in_3')
// (7, 11, 'lutff_2/in_0')
// (7, 11, 'lutff_3/in_2')
// (7, 11, 'lutff_4/in_0')
// (7, 11, 'lutff_6/in_0')
// (7, 11, 'sp12_h_r_6')
// (8, 10, 'neigh_op_tnr_1')
// (8, 11, 'local_g2_1')
// (8, 11, 'lutff_6/in_3')
// (8, 11, 'lutff_7/in_2')
// (8, 11, 'neigh_op_rgt_1')
// (8, 11, 'sp12_h_r_9')
// (8, 12, 'neigh_op_bnr_1')
// (9, 10, 'neigh_op_top_1')
// (9, 11, 'lutff_1/out')
// (9, 11, 'sp12_h_r_10')
// (9, 12, 'neigh_op_bot_1')
// (10, 10, 'neigh_op_tnl_1')
// (10, 11, 'neigh_op_lft_1')
// (10, 11, 'sp12_h_r_13')
// (10, 12, 'neigh_op_bnl_1')
// (11, 11, 'sp12_h_r_14')
// (12, 11, 'sp12_h_r_17')
// (13, 11, 'span12_horz_17')

wire n202;
// (4, 11, 'sp4_h_r_6')
// (5, 9, 'sp4_r_v_b_39')
// (5, 10, 'local_g0_2')
// (5, 10, 'lutff_5/in_1')
// (5, 10, 'sp4_r_v_b_26')
// (5, 11, 'local_g1_3')
// (5, 11, 'lutff_6/in_2')
// (5, 11, 'sp4_h_r_19')
// (5, 11, 'sp4_r_v_b_15')
// (5, 12, 'sp4_r_v_b_2')
// (6, 8, 'sp4_v_t_39')
// (6, 9, 'sp4_r_v_b_41')
// (6, 9, 'sp4_v_b_39')
// (6, 10, 'local_g0_4')
// (6, 10, 'lutff_5/in_1')
// (6, 10, 'sp4_r_v_b_28')
// (6, 10, 'sp4_v_b_26')
// (6, 11, 'neigh_op_tnr_2')
// (6, 11, 'sp4_h_r_30')
// (6, 11, 'sp4_r_v_b_17')
// (6, 11, 'sp4_v_b_15')
// (6, 12, 'neigh_op_rgt_2')
// (6, 12, 'sp4_h_r_9')
// (6, 12, 'sp4_r_v_b_4')
// (6, 12, 'sp4_v_b_2')
// (6, 13, 'neigh_op_bnr_2')
// (7, 8, 'sp4_v_t_41')
// (7, 9, 'sp4_v_b_41')
// (7, 10, 'sp4_v_b_28')
// (7, 11, 'neigh_op_top_2')
// (7, 11, 'sp4_h_r_43')
// (7, 11, 'sp4_v_b_17')
// (7, 12, 'lutff_2/out')
// (7, 12, 'sp4_h_r_20')
// (7, 12, 'sp4_r_v_b_37')
// (7, 12, 'sp4_v_b_4')
// (7, 13, 'neigh_op_bot_2')
// (7, 13, 'sp4_r_v_b_24')
// (7, 14, 'sp4_r_v_b_13')
// (7, 15, 'sp4_r_v_b_0')
// (8, 11, 'neigh_op_tnl_2')
// (8, 11, 'sp4_h_l_43')
// (8, 11, 'sp4_v_t_37')
// (8, 12, 'neigh_op_lft_2')
// (8, 12, 'sp4_h_r_33')
// (8, 12, 'sp4_v_b_37')
// (8, 13, 'neigh_op_bnl_2')
// (8, 13, 'sp4_v_b_24')
// (8, 14, 'sp4_v_b_13')
// (8, 15, 'sp4_v_b_0')
// (9, 12, 'sp4_h_r_44')
// (10, 12, 'sp4_h_l_44')

wire n203;
// (4, 12, 'sp12_h_r_1')
// (5, 12, 'sp12_h_r_2')
// (6, 12, 'sp12_h_r_5')
// (7, 12, 'sp12_h_r_6')
// (8, 11, 'neigh_op_tnr_1')
// (8, 12, 'neigh_op_rgt_1')
// (8, 12, 'sp12_h_r_9')
// (8, 13, 'neigh_op_bnr_1')
// (9, 11, 'neigh_op_top_1')
// (9, 12, 'lutff_1/out')
// (9, 12, 'sp12_h_r_10')
// (9, 13, 'neigh_op_bot_1')
// (10, 11, 'neigh_op_tnl_1')
// (10, 12, 'neigh_op_lft_1')
// (10, 12, 'sp12_h_r_13')
// (10, 13, 'neigh_op_bnl_1')
// (11, 12, 'local_g1_6')
// (11, 12, 'lutff_5/in_2')
// (11, 12, 'sp12_h_r_14')
// (12, 12, 'sp12_h_r_17')
// (13, 12, 'span12_horz_17')

wire n204;
// (4, 12, 'sp4_h_r_7')
// (5, 12, 'local_g1_2')
// (5, 12, 'lutff_5/in_2')
// (5, 12, 'sp4_h_r_18')
// (6, 11, 'neigh_op_tnr_5')
// (6, 12, 'neigh_op_rgt_5')
// (6, 12, 'sp4_h_r_31')
// (6, 13, 'neigh_op_bnr_5')
// (7, 11, 'neigh_op_top_5')
// (7, 12, 'lutff_5/out')
// (7, 12, 'sp4_h_r_42')
// (7, 13, 'neigh_op_bot_5')
// (8, 11, 'neigh_op_tnl_5')
// (8, 12, 'neigh_op_lft_5')
// (8, 12, 'sp4_h_l_42')
// (8, 13, 'neigh_op_bnl_5')

reg n205 = 0;
// (4, 14, 'local_g2_7')
// (4, 14, 'lutff_5/in_0')
// (4, 14, 'neigh_op_tnr_7')
// (4, 15, 'local_g2_7')
// (4, 15, 'lutff_0/in_1')
// (4, 15, 'neigh_op_rgt_7')
// (4, 16, 'neigh_op_bnr_7')
// (5, 14, 'local_g1_7')
// (5, 14, 'lutff_7/in_3')
// (5, 14, 'neigh_op_top_7')
// (5, 15, 'local_g0_7')
// (5, 15, 'local_g1_7')
// (5, 15, 'lutff_0/in_3')
// (5, 15, 'lutff_7/in_1')
// (5, 15, 'lutff_7/out')
// (5, 16, 'neigh_op_bot_7')
// (6, 14, 'neigh_op_tnl_7')
// (6, 15, 'neigh_op_lft_7')
// (6, 16, 'neigh_op_bnl_7')

wire n206;
// (4, 14, 'lutff_1/cout')
// (4, 14, 'lutff_2/in_3')

wire n207;
// (4, 14, 'lutff_2/cout')
// (4, 14, 'lutff_3/in_3')

wire n208;
// (4, 15, 'sp4_h_r_10')
// (5, 14, 'neigh_op_tnr_1')
// (5, 15, 'neigh_op_rgt_1')
// (5, 15, 'sp4_h_r_23')
// (5, 16, 'neigh_op_bnr_1')
// (6, 14, 'neigh_op_top_1')
// (6, 15, 'lutff_1/out')
// (6, 15, 'sp4_h_r_34')
// (6, 16, 'neigh_op_bot_1')
// (7, 12, 'sp4_r_v_b_47')
// (7, 13, 'sp4_r_v_b_34')
// (7, 14, 'local_g2_1')
// (7, 14, 'local_g3_1')
// (7, 14, 'lutff_1/in_2')
// (7, 14, 'lutff_2/in_2')
// (7, 14, 'lutff_6/in_0')
// (7, 14, 'lutff_7/in_3')
// (7, 14, 'neigh_op_tnl_1')
// (7, 14, 'sp4_r_v_b_23')
// (7, 15, 'neigh_op_lft_1')
// (7, 15, 'sp4_h_r_47')
// (7, 15, 'sp4_r_v_b_10')
// (7, 16, 'neigh_op_bnl_1')
// (8, 11, 'sp4_v_t_47')
// (8, 12, 'sp4_v_b_47')
// (8, 13, 'sp4_v_b_34')
// (8, 14, 'local_g0_7')
// (8, 14, 'local_g1_7')
// (8, 14, 'lutff_0/in_2')
// (8, 14, 'lutff_1/in_0')
// (8, 14, 'lutff_2/in_0')
// (8, 14, 'sp4_v_b_23')
// (8, 15, 'sp4_h_l_47')
// (8, 15, 'sp4_v_b_10')

wire n209;
// (5, 0, 'span12_vert_17')
// (5, 1, 'sp12_v_b_17')
// (5, 2, 'sp12_v_b_14')
// (5, 3, 'sp12_v_b_13')
// (5, 4, 'sp12_v_b_10')
// (5, 5, 'sp12_v_b_9')
// (5, 6, 'local_g2_6')
// (5, 6, 'local_g3_6')
// (5, 6, 'lutff_1/in_3')
// (5, 6, 'lutff_5/in_2')
// (5, 6, 'lutff_6/in_3')
// (5, 6, 'sp12_v_b_6')
// (5, 7, 'sp12_v_b_5')
// (5, 8, 'sp12_v_b_2')
// (5, 9, 'sp12_h_r_1')
// (5, 9, 'sp12_v_b_1')
// (6, 9, 'sp12_h_r_2')
// (7, 4, 'sp4_r_v_b_46')
// (7, 5, 'sp4_r_v_b_35')
// (7, 6, 'sp4_r_v_b_22')
// (7, 7, 'sp4_r_v_b_11')
// (7, 8, 'neigh_op_tnr_7')
// (7, 9, 'neigh_op_rgt_7')
// (7, 9, 'sp12_h_r_5')
// (7, 10, 'neigh_op_bnr_7')
// (8, 3, 'sp4_h_r_4')
// (8, 3, 'sp4_v_t_46')
// (8, 4, 'sp12_v_t_22')
// (8, 4, 'sp4_v_b_46')
// (8, 5, 'sp12_v_b_22')
// (8, 5, 'sp4_v_b_35')
// (8, 6, 'sp12_v_b_21')
// (8, 6, 'sp4_v_b_22')
// (8, 7, 'sp12_v_b_18')
// (8, 7, 'sp4_v_b_11')
// (8, 8, 'neigh_op_top_7')
// (8, 8, 'sp12_v_b_17')
// (8, 9, 'lutff_7/out')
// (8, 9, 'sp12_h_r_6')
// (8, 9, 'sp12_v_b_14')
// (8, 10, 'neigh_op_bot_7')
// (8, 10, 'sp12_v_b_13')
// (8, 11, 'sp12_v_b_10')
// (8, 12, 'sp12_v_b_9')
// (8, 13, 'sp12_v_b_6')
// (8, 14, 'sp12_v_b_5')
// (8, 15, 'sp12_v_b_2')
// (8, 16, 'sp12_v_b_1')
// (9, 3, 'sp4_h_r_17')
// (9, 8, 'neigh_op_tnl_7')
// (9, 9, 'neigh_op_lft_7')
// (9, 9, 'sp12_h_r_9')
// (9, 10, 'neigh_op_bnl_7')
// (10, 3, 'sp4_h_r_28')
// (10, 9, 'sp12_h_r_10')
// (11, 3, 'local_g2_1')
// (11, 3, 'lutff_1/in_2')
// (11, 3, 'sp4_h_r_41')
// (11, 9, 'local_g1_5')
// (11, 9, 'lutff_6/in_2')
// (11, 9, 'lutff_7/in_3')
// (11, 9, 'sp12_h_r_13')
// (12, 3, 'sp4_h_l_41')
// (12, 9, 'sp12_h_r_14')
// (13, 9, 'span12_horz_14')

reg n210 = 0;
// (5, 1, 'neigh_op_tnr_7')
// (5, 2, 'neigh_op_rgt_7')
// (5, 3, 'neigh_op_bnr_7')
// (6, 1, 'neigh_op_top_7')
// (6, 1, 'sp4_r_v_b_26')
// (6, 2, 'lutff_7/out')
// (6, 2, 'sp4_r_v_b_15')
// (6, 3, 'local_g1_2')
// (6, 3, 'lutff_2/in_1')
// (6, 3, 'neigh_op_bot_7')
// (6, 3, 'sp4_r_v_b_2')
// (7, 0, 'span4_vert_26')
// (7, 1, 'neigh_op_tnl_7')
// (7, 1, 'sp4_v_b_26')
// (7, 2, 'neigh_op_lft_7')
// (7, 2, 'sp4_v_b_15')
// (7, 3, 'neigh_op_bnl_7')
// (7, 3, 'sp4_v_b_2')

reg n211 = 0;
// (5, 2, 'neigh_op_tnr_1')
// (5, 3, 'neigh_op_rgt_1')
// (5, 4, 'neigh_op_bnr_1')
// (6, 2, 'neigh_op_top_1')
// (6, 3, 'local_g0_1')
// (6, 3, 'lutff_0/in_1')
// (6, 3, 'lutff_1/out')
// (6, 4, 'neigh_op_bot_1')
// (7, 2, 'neigh_op_tnl_1')
// (7, 3, 'neigh_op_lft_1')
// (7, 4, 'neigh_op_bnl_1')

reg n212 = 0;
// (5, 2, 'neigh_op_tnr_2')
// (5, 3, 'neigh_op_rgt_2')
// (5, 4, 'neigh_op_bnr_2')
// (6, 2, 'neigh_op_top_2')
// (6, 3, 'local_g0_2')
// (6, 3, 'lutff_1/in_1')
// (6, 3, 'lutff_2/out')
// (6, 4, 'neigh_op_bot_2')
// (7, 2, 'neigh_op_tnl_2')
// (7, 3, 'neigh_op_lft_2')
// (7, 4, 'neigh_op_bnl_2')

reg n213 = 0;
// (5, 2, 'neigh_op_tnr_3')
// (5, 3, 'neigh_op_rgt_3')
// (5, 4, 'neigh_op_bnr_3')
// (6, 2, 'neigh_op_top_3')
// (6, 3, 'local_g0_3')
// (6, 3, 'local_g1_3')
// (6, 3, 'lutff_1/in_2')
// (6, 3, 'lutff_3/out')
// (6, 3, 'lutff_7/in_1')
// (6, 4, 'neigh_op_bot_3')
// (7, 2, 'neigh_op_tnl_3')
// (7, 3, 'neigh_op_lft_3')
// (7, 4, 'neigh_op_bnl_3')

reg n214 = 0;
// (5, 2, 'neigh_op_tnr_4')
// (5, 3, 'neigh_op_rgt_4')
// (5, 4, 'neigh_op_bnr_4')
// (6, 2, 'local_g1_4')
// (6, 2, 'lutff_7/in_0')
// (6, 2, 'neigh_op_top_4')
// (6, 3, 'local_g0_4')
// (6, 3, 'lutff_4/out')
// (6, 3, 'lutff_5/in_1')
// (6, 4, 'neigh_op_bot_4')
// (7, 2, 'neigh_op_tnl_4')
// (7, 3, 'neigh_op_lft_4')
// (7, 4, 'neigh_op_bnl_4')

reg n215 = 0;
// (5, 2, 'neigh_op_tnr_5')
// (5, 3, 'neigh_op_rgt_5')
// (5, 4, 'neigh_op_bnr_5')
// (6, 2, 'neigh_op_top_5')
// (6, 3, 'local_g1_5')
// (6, 3, 'lutff_2/in_2')
// (6, 3, 'lutff_3/in_1')
// (6, 3, 'lutff_5/out')
// (6, 4, 'neigh_op_bot_5')
// (7, 2, 'neigh_op_tnl_5')
// (7, 3, 'neigh_op_lft_5')
// (7, 4, 'neigh_op_bnl_5')

reg n216 = 0;
// (5, 2, 'neigh_op_tnr_7')
// (5, 3, 'neigh_op_rgt_7')
// (5, 4, 'neigh_op_bnr_7')
// (6, 2, 'neigh_op_top_7')
// (6, 3, 'local_g0_7')
// (6, 3, 'local_g1_7')
// (6, 3, 'lutff_0/in_0')
// (6, 3, 'lutff_4/in_1')
// (6, 3, 'lutff_7/out')
// (6, 4, 'neigh_op_bot_7')
// (7, 2, 'neigh_op_tnl_7')
// (7, 3, 'neigh_op_lft_7')
// (7, 4, 'neigh_op_bnl_7')

reg n217 = 0;
// (5, 3, 'neigh_op_tnr_0')
// (5, 4, 'neigh_op_rgt_0')
// (5, 5, 'neigh_op_bnr_0')
// (6, 3, 'neigh_op_top_0')
// (6, 4, 'lutff_0/out')
// (6, 5, 'local_g0_0')
// (6, 5, 'lutff_0/in_0')
// (6, 5, 'neigh_op_bot_0')
// (7, 3, 'neigh_op_tnl_0')
// (7, 4, 'neigh_op_lft_0')
// (7, 5, 'neigh_op_bnl_0')

reg n218 = 0;
// (5, 3, 'neigh_op_tnr_2')
// (5, 4, 'neigh_op_rgt_2')
// (5, 5, 'neigh_op_bnr_2')
// (6, 3, 'neigh_op_top_2')
// (6, 4, 'local_g0_2')
// (6, 4, 'lutff_2/out')
// (6, 4, 'lutff_4/in_0')
// (6, 5, 'neigh_op_bot_2')
// (7, 3, 'neigh_op_tnl_2')
// (7, 4, 'neigh_op_lft_2')
// (7, 5, 'neigh_op_bnl_2')

reg n219 = 0;
// (5, 3, 'neigh_op_tnr_4')
// (5, 4, 'neigh_op_rgt_4')
// (5, 5, 'neigh_op_bnr_4')
// (6, 3, 'neigh_op_top_4')
// (6, 4, 'local_g1_4')
// (6, 4, 'lutff_3/in_0')
// (6, 4, 'lutff_4/out')
// (6, 5, 'neigh_op_bot_4')
// (7, 3, 'neigh_op_tnl_4')
// (7, 4, 'neigh_op_lft_4')
// (7, 5, 'neigh_op_bnl_4')

reg \d_out[3] = 0 ;
// (5, 3, 'neigh_op_tnr_7')
// (5, 4, 'neigh_op_rgt_7')
// (5, 5, 'neigh_op_bnr_7')
// (6, 1, 'sp4_r_v_b_25')
// (6, 2, 'sp4_r_v_b_12')
// (6, 3, 'neigh_op_top_7')
// (6, 3, 'sp4_r_v_b_1')
// (6, 4, 'lutff_7/out')
// (6, 4, 'sp4_r_v_b_47')
// (6, 5, 'neigh_op_bot_7')
// (6, 5, 'sp4_r_v_b_34')
// (6, 6, 'sp4_r_v_b_23')
// (6, 7, 'sp4_r_v_b_10')
// (7, 0, 'io_1/D_OUT_0')
// (7, 0, 'io_1/PAD')
// (7, 0, 'local_g0_1')
// (7, 0, 'span4_vert_25')
// (7, 1, 'sp4_v_b_25')
// (7, 2, 'sp4_v_b_12')
// (7, 3, 'neigh_op_tnl_7')
// (7, 3, 'sp4_v_b_1')
// (7, 3, 'sp4_v_t_47')
// (7, 4, 'neigh_op_lft_7')
// (7, 4, 'sp4_v_b_47')
// (7, 5, 'neigh_op_bnl_7')
// (7, 5, 'sp4_v_b_34')
// (7, 6, 'sp4_v_b_23')
// (7, 7, 'sp4_v_b_10')

reg n221 = 0;
// (5, 4, 'neigh_op_tnr_0')
// (5, 5, 'neigh_op_rgt_0')
// (5, 6, 'neigh_op_bnr_0')
// (6, 4, 'neigh_op_top_0')
// (6, 5, 'lutff_0/out')
// (6, 6, 'local_g1_0')
// (6, 6, 'lutff_5/in_0')
// (6, 6, 'neigh_op_bot_0')
// (7, 4, 'neigh_op_tnl_0')
// (7, 5, 'neigh_op_lft_0')
// (7, 6, 'neigh_op_bnl_0')

reg n222 = 0;
// (5, 4, 'neigh_op_tnr_1')
// (5, 5, 'neigh_op_rgt_1')
// (5, 6, 'neigh_op_bnr_1')
// (6, 4, 'neigh_op_top_1')
// (6, 5, 'local_g0_1')
// (6, 5, 'lutff_1/out')
// (6, 5, 'lutff_7/in_0')
// (6, 6, 'neigh_op_bot_1')
// (7, 4, 'neigh_op_tnl_1')
// (7, 5, 'neigh_op_lft_1')
// (7, 6, 'neigh_op_bnl_1')

reg n223 = 0;
// (5, 4, 'neigh_op_tnr_2')
// (5, 5, 'neigh_op_rgt_2')
// (5, 6, 'neigh_op_bnr_2')
// (6, 4, 'neigh_op_top_2')
// (6, 5, 'local_g1_2')
// (6, 5, 'lutff_2/out')
// (6, 5, 'lutff_5/in_0')
// (6, 6, 'neigh_op_bot_2')
// (7, 4, 'neigh_op_tnl_2')
// (7, 5, 'neigh_op_lft_2')
// (7, 6, 'neigh_op_bnl_2')

reg n224 = 0;
// (5, 4, 'neigh_op_tnr_3')
// (5, 5, 'neigh_op_rgt_3')
// (5, 6, 'neigh_op_bnr_3')
// (6, 4, 'neigh_op_top_3')
// (6, 5, 'local_g1_3')
// (6, 5, 'lutff_3/out')
// (6, 5, 'lutff_6/in_0')
// (6, 6, 'neigh_op_bot_3')
// (7, 4, 'neigh_op_tnl_3')
// (7, 5, 'neigh_op_lft_3')
// (7, 6, 'neigh_op_bnl_3')

reg n225 = 0;
// (5, 4, 'neigh_op_tnr_4')
// (5, 5, 'neigh_op_rgt_4')
// (5, 6, 'neigh_op_bnr_4')
// (6, 4, 'neigh_op_top_4')
// (6, 5, 'local_g0_4')
// (6, 5, 'lutff_3/in_1')
// (6, 5, 'lutff_4/out')
// (6, 6, 'neigh_op_bot_4')
// (7, 4, 'neigh_op_tnl_4')
// (7, 5, 'local_g1_4')
// (7, 5, 'lutff_0/in_1')
// (7, 5, 'neigh_op_lft_4')
// (7, 6, 'neigh_op_bnl_4')

reg n226 = 0;
// (5, 4, 'neigh_op_tnr_5')
// (5, 5, 'neigh_op_rgt_5')
// (5, 6, 'neigh_op_bnr_5')
// (6, 2, 'sp4_r_v_b_46')
// (6, 3, 'sp4_r_v_b_35')
// (6, 4, 'neigh_op_top_5')
// (6, 4, 'sp4_r_v_b_22')
// (6, 5, 'local_g0_5')
// (6, 5, 'lutff_3/in_0')
// (6, 5, 'lutff_5/out')
// (6, 5, 'sp4_r_v_b_11')
// (6, 6, 'neigh_op_bot_5')
// (7, 1, 'sp4_v_t_46')
// (7, 2, 'sp4_v_b_46')
// (7, 3, 'sp4_v_b_35')
// (7, 4, 'neigh_op_tnl_5')
// (7, 4, 'sp4_v_b_22')
// (7, 5, 'local_g1_3')
// (7, 5, 'lutff_1/in_1')
// (7, 5, 'lutff_2/in_0')
// (7, 5, 'lutff_6/in_2')
// (7, 5, 'neigh_op_lft_5')
// (7, 5, 'sp4_v_b_11')
// (7, 6, 'neigh_op_bnl_5')

reg n227 = 0;
// (5, 4, 'neigh_op_tnr_6')
// (5, 5, 'neigh_op_rgt_6')
// (5, 6, 'neigh_op_bnr_6')
// (6, 4, 'neigh_op_top_6')
// (6, 5, 'local_g0_6')
// (6, 5, 'lutff_2/in_0')
// (6, 5, 'lutff_6/out')
// (6, 6, 'neigh_op_bot_6')
// (7, 4, 'neigh_op_tnl_6')
// (7, 5, 'neigh_op_lft_6')
// (7, 6, 'neigh_op_bnl_6')

reg n228 = 0;
// (5, 4, 'neigh_op_tnr_7')
// (5, 5, 'neigh_op_rgt_7')
// (5, 6, 'neigh_op_bnr_7')
// (6, 4, 'neigh_op_top_7')
// (6, 5, 'local_g1_7')
// (6, 5, 'lutff_4/in_0')
// (6, 5, 'lutff_7/out')
// (6, 6, 'neigh_op_bot_7')
// (7, 4, 'neigh_op_tnl_7')
// (7, 5, 'neigh_op_lft_7')
// (7, 6, 'neigh_op_bnl_7')

wire n229;
// (5, 5, 'neigh_op_tnr_1')
// (5, 6, 'neigh_op_rgt_1')
// (5, 7, 'neigh_op_bnr_1')
// (6, 5, 'neigh_op_top_1')
// (6, 6, 'lutff_1/out')
// (6, 7, 'neigh_op_bot_1')
// (7, 5, 'local_g2_1')
// (7, 5, 'local_g3_1')
// (7, 5, 'lutff_0/in_0')
// (7, 5, 'lutff_6/in_1')
// (7, 5, 'neigh_op_tnl_1')
// (7, 6, 'neigh_op_lft_1')
// (7, 7, 'neigh_op_bnl_1')

reg n230 = 0;
// (5, 5, 'neigh_op_tnr_2')
// (5, 6, 'neigh_op_rgt_2')
// (5, 7, 'neigh_op_bnr_2')
// (6, 5, 'neigh_op_top_2')
// (6, 6, 'lutff_2/out')
// (6, 6, 'sp4_h_r_4')
// (6, 7, 'neigh_op_bot_2')
// (7, 5, 'neigh_op_tnl_2')
// (7, 6, 'local_g1_1')
// (7, 6, 'lutff_6/in_0')
// (7, 6, 'neigh_op_lft_2')
// (7, 6, 'sp4_h_r_17')
// (7, 7, 'neigh_op_bnl_2')
// (8, 6, 'sp4_h_r_28')
// (9, 6, 'sp4_h_r_41')
// (10, 6, 'sp4_h_l_41')

reg n231 = 0;
// (5, 5, 'neigh_op_tnr_4')
// (5, 6, 'neigh_op_rgt_4')
// (5, 7, 'neigh_op_bnr_4')
// (6, 5, 'neigh_op_top_4')
// (6, 6, 'local_g0_4')
// (6, 6, 'lutff_4/out')
// (6, 6, 'lutff_6/in_0')
// (6, 7, 'neigh_op_bot_4')
// (7, 5, 'neigh_op_tnl_4')
// (7, 6, 'neigh_op_lft_4')
// (7, 7, 'neigh_op_bnl_4')

reg n232 = 0;
// (5, 5, 'neigh_op_tnr_5')
// (5, 5, 'sp4_r_v_b_39')
// (5, 6, 'neigh_op_rgt_5')
// (5, 6, 'sp4_r_v_b_26')
// (5, 7, 'neigh_op_bnr_5')
// (5, 7, 'sp4_r_v_b_15')
// (5, 8, 'sp4_r_v_b_2')
// (5, 9, 'sp4_r_v_b_40')
// (5, 10, 'sp4_r_v_b_29')
// (5, 11, 'sp4_r_v_b_16')
// (5, 12, 'sp4_r_v_b_5')
// (6, 4, 'sp4_v_t_39')
// (6, 5, 'neigh_op_top_5')
// (6, 5, 'sp4_v_b_39')
// (6, 6, 'lutff_5/out')
// (6, 6, 'sp4_v_b_26')
// (6, 7, 'neigh_op_bot_5')
// (6, 7, 'sp4_v_b_15')
// (6, 8, 'sp4_v_b_2')
// (6, 8, 'sp4_v_t_40')
// (6, 9, 'sp4_v_b_40')
// (6, 10, 'sp4_v_b_29')
// (6, 11, 'sp4_v_b_16')
// (6, 12, 'local_g1_5')
// (6, 12, 'lutff_3/in_3')
// (6, 12, 'sp4_v_b_5')
// (7, 5, 'neigh_op_tnl_5')
// (7, 6, 'neigh_op_lft_5')
// (7, 7, 'neigh_op_bnl_5')

reg n233 = 0;
// (5, 5, 'neigh_op_tnr_6')
// (5, 6, 'neigh_op_rgt_6')
// (5, 7, 'neigh_op_bnr_6')
// (6, 5, 'neigh_op_top_6')
// (6, 6, 'local_g0_6')
// (6, 6, 'lutff_2/in_0')
// (6, 6, 'lutff_6/out')
// (6, 7, 'neigh_op_bot_6')
// (7, 5, 'neigh_op_tnl_6')
// (7, 6, 'neigh_op_lft_6')
// (7, 7, 'neigh_op_bnl_6')

wire n234;
// (5, 6, 'neigh_op_tnr_0')
// (5, 7, 'neigh_op_rgt_0')
// (5, 8, 'neigh_op_bnr_0')
// (6, 6, 'neigh_op_top_0')
// (6, 6, 'sp4_r_v_b_44')
// (6, 7, 'lutff_0/out')
// (6, 7, 'sp4_r_v_b_33')
// (6, 8, 'neigh_op_bot_0')
// (6, 8, 'sp4_r_v_b_20')
// (6, 9, 'sp4_r_v_b_9')
// (7, 5, 'sp4_v_t_44')
// (7, 6, 'neigh_op_tnl_0')
// (7, 6, 'sp4_v_b_44')
// (7, 7, 'neigh_op_lft_0')
// (7, 7, 'sp4_v_b_33')
// (7, 8, 'neigh_op_bnl_0')
// (7, 8, 'sp4_v_b_20')
// (7, 9, 'local_g1_3')
// (7, 9, 'lutff_6/in_0')
// (7, 9, 'sp4_h_r_3')
// (7, 9, 'sp4_v_b_9')
// (8, 9, 'sp4_h_r_14')
// (9, 9, 'sp4_h_r_27')
// (10, 9, 'sp4_h_r_38')
// (11, 9, 'sp4_h_l_38')

wire n235;
// (5, 6, 'neigh_op_tnr_1')
// (5, 7, 'neigh_op_rgt_1')
// (5, 8, 'neigh_op_bnr_1')
// (6, 6, 'neigh_op_top_1')
// (6, 7, 'local_g2_1')
// (6, 7, 'lutff_0/in_3')
// (6, 7, 'lutff_1/out')
// (6, 8, 'neigh_op_bot_1')
// (7, 6, 'neigh_op_tnl_1')
// (7, 7, 'neigh_op_lft_1')
// (7, 8, 'neigh_op_bnl_1')

reg n236 = 0;
// (5, 6, 'neigh_op_tnr_3')
// (5, 7, 'local_g2_3')
// (5, 7, 'lutff_1/in_0')
// (5, 7, 'neigh_op_rgt_3')
// (5, 8, 'neigh_op_bnr_3')
// (6, 6, 'neigh_op_top_3')
// (6, 7, 'lutff_3/out')
// (6, 8, 'neigh_op_bot_3')
// (7, 6, 'neigh_op_tnl_3')
// (7, 7, 'neigh_op_lft_3')
// (7, 8, 'neigh_op_bnl_3')

reg n237 = 0;
// (5, 6, 'neigh_op_tnr_4')
// (5, 7, 'neigh_op_rgt_4')
// (5, 8, 'neigh_op_bnr_4')
// (6, 6, 'neigh_op_top_4')
// (6, 7, 'local_g0_4')
// (6, 7, 'lutff_4/out')
// (6, 7, 'lutff_6/in_0')
// (6, 8, 'neigh_op_bot_4')
// (7, 6, 'neigh_op_tnl_4')
// (7, 7, 'neigh_op_lft_4')
// (7, 8, 'neigh_op_bnl_4')

reg n238 = 0;
// (5, 6, 'neigh_op_tnr_5')
// (5, 7, 'neigh_op_rgt_5')
// (5, 8, 'neigh_op_bnr_5')
// (6, 6, 'neigh_op_top_5')
// (6, 7, 'local_g0_5')
// (6, 7, 'lutff_5/out')
// (6, 7, 'lutff_7/in_0')
// (6, 8, 'neigh_op_bot_5')
// (7, 6, 'neigh_op_tnl_5')
// (7, 7, 'neigh_op_lft_5')
// (7, 8, 'neigh_op_bnl_5')

reg n239 = 0;
// (5, 6, 'neigh_op_tnr_6')
// (5, 7, 'neigh_op_rgt_6')
// (5, 8, 'neigh_op_bnr_6')
// (6, 6, 'neigh_op_top_6')
// (6, 7, 'local_g1_6')
// (6, 7, 'lutff_5/in_0')
// (6, 7, 'lutff_6/out')
// (6, 8, 'neigh_op_bot_6')
// (7, 6, 'neigh_op_tnl_6')
// (7, 7, 'neigh_op_lft_6')
// (7, 8, 'neigh_op_bnl_6')

reg n240 = 0;
// (5, 6, 'neigh_op_tnr_7')
// (5, 7, 'neigh_op_rgt_7')
// (5, 8, 'neigh_op_bnr_7')
// (6, 6, 'neigh_op_top_7')
// (6, 7, 'local_g2_7')
// (6, 7, 'local_g3_7')
// (6, 7, 'lutff_1/in_0')
// (6, 7, 'lutff_3/in_1')
// (6, 7, 'lutff_7/out')
// (6, 8, 'neigh_op_bot_7')
// (7, 6, 'neigh_op_tnl_7')
// (7, 7, 'neigh_op_lft_7')
// (7, 8, 'neigh_op_bnl_7')

reg n241 = 0;
// (5, 6, 'sp4_h_r_2')
// (6, 5, 'neigh_op_tnr_5')
// (6, 6, 'neigh_op_rgt_5')
// (6, 6, 'sp4_h_r_15')
// (6, 7, 'neigh_op_bnr_5')
// (7, 5, 'neigh_op_top_5')
// (7, 6, 'lutff_5/out')
// (7, 6, 'sp4_h_r_26')
// (7, 7, 'neigh_op_bot_5')
// (8, 5, 'neigh_op_tnl_5')
// (8, 6, 'local_g2_7')
// (8, 6, 'lutff_6/in_3')
// (8, 6, 'neigh_op_lft_5')
// (8, 6, 'sp4_h_r_39')
// (8, 7, 'neigh_op_bnl_5')
// (9, 6, 'sp4_h_l_39')

wire n242;
// (5, 6, 'sp4_r_v_b_41')
// (5, 7, 'local_g1_4')
// (5, 7, 'lutff_2/in_3')
// (5, 7, 'lutff_4/in_3')
// (5, 7, 'sp4_r_v_b_28')
// (5, 8, 'sp4_r_v_b_17')
// (5, 9, 'sp4_r_v_b_4')
// (5, 10, 'local_g2_5')
// (5, 10, 'lutff_5/in_2')
// (5, 10, 'sp4_r_v_b_37')
// (5, 11, 'sp4_r_v_b_24')
// (5, 12, 'sp4_r_v_b_13')
// (5, 13, 'sp4_r_v_b_0')
// (6, 5, 'sp4_v_t_41')
// (6, 6, 'sp4_v_b_41')
// (6, 7, 'sp4_v_b_28')
// (6, 8, 'local_g2_3')
// (6, 8, 'lutff_7/in_2')
// (6, 8, 'neigh_op_tnr_3')
// (6, 8, 'sp4_v_b_17')
// (6, 9, 'local_g2_3')
// (6, 9, 'lutff_2/in_3')
// (6, 9, 'lutff_5/in_2')
// (6, 9, 'neigh_op_rgt_3')
// (6, 9, 'sp4_h_r_11')
// (6, 9, 'sp4_v_b_4')
// (6, 9, 'sp4_v_t_37')
// (6, 10, 'neigh_op_bnr_3')
// (6, 10, 'sp4_v_b_37')
// (6, 11, 'sp4_v_b_24')
// (6, 12, 'sp4_v_b_13')
// (6, 13, 'sp4_v_b_0')
// (7, 8, 'neigh_op_top_3')
// (7, 9, 'lutff_3/out')
// (7, 9, 'sp4_h_r_22')
// (7, 10, 'neigh_op_bot_3')
// (8, 8, 'neigh_op_tnl_3')
// (8, 9, 'neigh_op_lft_3')
// (8, 9, 'sp4_h_r_35')
// (8, 10, 'neigh_op_bnl_3')
// (9, 9, 'sp4_h_r_46')
// (10, 9, 'sp4_h_l_46')

reg n243 = 0;
// (5, 6, 'sp4_r_v_b_43')
// (5, 7, 'sp4_r_v_b_30')
// (5, 8, 'neigh_op_tnr_3')
// (5, 8, 'sp4_r_v_b_19')
// (5, 9, 'neigh_op_rgt_3')
// (5, 9, 'sp4_r_v_b_6')
// (5, 10, 'neigh_op_bnr_3')
// (6, 5, 'sp4_v_t_43')
// (6, 6, 'local_g2_3')
// (6, 6, 'lutff_1/in_0')
// (6, 6, 'sp4_v_b_43')
// (6, 7, 'sp4_v_b_30')
// (6, 8, 'neigh_op_top_3')
// (6, 8, 'sp4_v_b_19')
// (6, 9, 'local_g0_3')
// (6, 9, 'lutff_2/in_1')
// (6, 9, 'lutff_3/out')
// (6, 9, 'sp4_v_b_6')
// (6, 10, 'neigh_op_bot_3')
// (7, 8, 'neigh_op_tnl_3')
// (7, 9, 'neigh_op_lft_3')
// (7, 10, 'neigh_op_bnl_3')

reg n244 = 0;
// (5, 7, 'neigh_op_tnr_0')
// (5, 8, 'neigh_op_rgt_0')
// (5, 9, 'neigh_op_bnr_0')
// (6, 5, 'sp4_r_v_b_36')
// (6, 6, 'local_g1_1')
// (6, 6, 'lutff_4/in_0')
// (6, 6, 'sp4_r_v_b_25')
// (6, 7, 'neigh_op_top_0')
// (6, 7, 'sp4_r_v_b_12')
// (6, 8, 'lutff_0/out')
// (6, 8, 'sp4_r_v_b_1')
// (6, 9, 'neigh_op_bot_0')
// (7, 4, 'sp4_v_t_36')
// (7, 5, 'sp4_v_b_36')
// (7, 6, 'sp4_v_b_25')
// (7, 7, 'neigh_op_tnl_0')
// (7, 7, 'sp4_v_b_12')
// (7, 8, 'neigh_op_lft_0')
// (7, 8, 'sp4_v_b_1')
// (7, 9, 'neigh_op_bnl_0')

reg n245 = 0;
// (5, 7, 'neigh_op_tnr_1')
// (5, 8, 'neigh_op_rgt_1')
// (5, 9, 'neigh_op_bnr_1')
// (6, 7, 'neigh_op_top_1')
// (6, 8, 'local_g0_1')
// (6, 8, 'lutff_1/out')
// (6, 8, 'lutff_2/in_1')
// (6, 8, 'lutff_3/in_2')
// (6, 9, 'neigh_op_bot_1')
// (7, 7, 'neigh_op_tnl_1')
// (7, 8, 'neigh_op_lft_1')
// (7, 9, 'neigh_op_bnl_1')

reg n246 = 0;
// (5, 7, 'neigh_op_tnr_6')
// (5, 8, 'neigh_op_rgt_6')
// (5, 9, 'neigh_op_bnr_6')
// (6, 7, 'neigh_op_top_6')
// (6, 8, 'local_g0_6')
// (6, 8, 'lutff_3/in_1')
// (6, 8, 'lutff_6/out')
// (6, 9, 'neigh_op_bot_6')
// (7, 7, 'neigh_op_tnl_6')
// (7, 8, 'neigh_op_lft_6')
// (7, 9, 'neigh_op_bnl_6')

reg n247 = 0;
// (5, 7, 'neigh_op_tnr_7')
// (5, 8, 'neigh_op_rgt_7')
// (5, 9, 'neigh_op_bnr_7')
// (6, 7, 'neigh_op_top_7')
// (6, 8, 'local_g1_7')
// (6, 8, 'lutff_1/in_1')
// (6, 8, 'lutff_6/in_2')
// (6, 8, 'lutff_7/out')
// (6, 9, 'neigh_op_bot_7')
// (7, 7, 'neigh_op_tnl_7')
// (7, 8, 'neigh_op_lft_7')
// (7, 9, 'neigh_op_bnl_7')

reg n248 = 0;
// (5, 7, 'sp12_h_r_1')
// (6, 7, 'sp12_h_r_2')
// (7, 7, 'sp12_h_r_5')
// (8, 7, 'sp12_h_r_6')
// (9, 7, 'local_g0_3')
// (9, 7, 'local_g1_1')
// (9, 7, 'lutff_1/in_1')
// (9, 7, 'lutff_3/in_0')
// (9, 7, 'lutff_5/in_0')
// (9, 7, 'sp12_h_r_9')
// (9, 7, 'sp4_h_r_3')
// (10, 7, 'sp12_h_r_10')
// (10, 7, 'sp4_h_r_14')
// (11, 6, 'neigh_op_tnr_3')
// (11, 7, 'local_g3_3')
// (11, 7, 'lutff_4/in_2')
// (11, 7, 'neigh_op_rgt_3')
// (11, 7, 'sp12_h_r_13')
// (11, 7, 'sp4_h_r_27')
// (11, 8, 'neigh_op_bnr_3')
// (12, 6, 'neigh_op_top_3')
// (12, 7, 'lutff_3/out')
// (12, 7, 'sp12_h_r_14')
// (12, 7, 'sp4_h_r_38')
// (12, 8, 'neigh_op_bot_3')
// (13, 6, 'logic_op_tnl_3')
// (13, 7, 'logic_op_lft_3')
// (13, 7, 'span12_horz_14')
// (13, 7, 'span4_horz_38')
// (13, 8, 'logic_op_bnl_3')

reg n249 = 0;
// (5, 8, 'neigh_op_tnr_0')
// (5, 9, 'neigh_op_rgt_0')
// (5, 10, 'neigh_op_bnr_0')
// (6, 8, 'neigh_op_top_0')
// (6, 9, 'local_g0_0')
// (6, 9, 'lutff_0/out')
// (6, 9, 'lutff_1/in_1')
// (6, 10, 'neigh_op_bot_0')
// (7, 8, 'neigh_op_tnl_0')
// (7, 9, 'neigh_op_lft_0')
// (7, 10, 'neigh_op_bnl_0')

reg n250 = 0;
// (5, 8, 'neigh_op_tnr_1')
// (5, 9, 'neigh_op_rgt_1')
// (5, 10, 'neigh_op_bnr_1')
// (6, 6, 'local_g2_6')
// (6, 6, 'lutff_1/in_1')
// (6, 6, 'sp4_r_v_b_38')
// (6, 7, 'sp4_r_v_b_27')
// (6, 8, 'neigh_op_top_1')
// (6, 8, 'sp4_r_v_b_14')
// (6, 9, 'lutff_1/out')
// (6, 9, 'sp4_r_v_b_3')
// (6, 10, 'neigh_op_bot_1')
// (7, 5, 'sp4_v_t_38')
// (7, 6, 'sp4_v_b_38')
// (7, 7, 'sp4_v_b_27')
// (7, 8, 'neigh_op_tnl_1')
// (7, 8, 'sp4_v_b_14')
// (7, 9, 'neigh_op_lft_1')
// (7, 9, 'sp4_v_b_3')
// (7, 10, 'neigh_op_bnl_1')

reg n251 = 0;
// (5, 8, 'neigh_op_tnr_4')
// (5, 9, 'neigh_op_rgt_4')
// (5, 10, 'neigh_op_bnr_4')
// (6, 8, 'neigh_op_top_4')
// (6, 9, 'local_g2_4')
// (6, 9, 'local_g3_4')
// (6, 9, 'lutff_1/in_2')
// (6, 9, 'lutff_3/in_1')
// (6, 9, 'lutff_4/out')
// (6, 10, 'neigh_op_bot_4')
// (7, 8, 'neigh_op_tnl_4')
// (7, 9, 'neigh_op_lft_4')
// (7, 10, 'neigh_op_bnl_4')

reg n252 = 0;
// (5, 8, 'neigh_op_tnr_5')
// (5, 9, 'neigh_op_rgt_5')
// (5, 10, 'neigh_op_bnr_5')
// (6, 8, 'neigh_op_top_5')
// (6, 9, 'local_g0_5')
// (6, 9, 'local_g1_5')
// (6, 9, 'lutff_0/in_2')
// (6, 9, 'lutff_4/in_1')
// (6, 9, 'lutff_5/out')
// (6, 10, 'neigh_op_bot_5')
// (7, 8, 'neigh_op_tnl_5')
// (7, 9, 'neigh_op_lft_5')
// (7, 10, 'neigh_op_bnl_5')

reg n253 = 0;
// (5, 8, 'neigh_op_tnr_6')
// (5, 9, 'neigh_op_rgt_6')
// (5, 10, 'neigh_op_bnr_6')
// (6, 8, 'neigh_op_top_6')
// (6, 9, 'local_g3_6')
// (6, 9, 'lutff_6/out')
// (6, 9, 'lutff_7/in_0')
// (6, 10, 'neigh_op_bot_6')
// (7, 8, 'neigh_op_tnl_6')
// (7, 9, 'neigh_op_lft_6')
// (7, 10, 'neigh_op_bnl_6')

reg n254 = 0;
// (5, 8, 'neigh_op_tnr_7')
// (5, 9, 'neigh_op_rgt_7')
// (5, 10, 'neigh_op_bnr_7')
// (6, 4, 'sp12_v_t_22')
// (6, 5, 'sp12_v_b_22')
// (6, 6, 'sp12_v_b_21')
// (6, 7, 'sp12_v_b_18')
// (6, 8, 'neigh_op_top_7')
// (6, 8, 'sp12_v_b_17')
// (6, 9, 'lutff_7/out')
// (6, 9, 'sp12_v_b_14')
// (6, 10, 'local_g1_7')
// (6, 10, 'lutff_0/in_0')
// (6, 10, 'neigh_op_bot_7')
// (6, 10, 'sp12_v_b_13')
// (6, 11, 'local_g3_2')
// (6, 11, 'lutff_6/in_3')
// (6, 11, 'sp12_v_b_10')
// (6, 12, 'sp12_v_b_9')
// (6, 13, 'sp12_v_b_6')
// (6, 14, 'sp12_v_b_5')
// (6, 15, 'sp12_v_b_2')
// (6, 16, 'sp12_v_b_1')
// (7, 8, 'neigh_op_tnl_7')
// (7, 9, 'neigh_op_lft_7')
// (7, 10, 'neigh_op_bnl_7')

reg n255 = 0;
// (5, 8, 'sp12_h_r_0')
// (6, 7, 'neigh_op_tnr_6')
// (6, 8, 'neigh_op_rgt_6')
// (6, 8, 'sp12_h_r_3')
// (6, 9, 'neigh_op_bnr_6')
// (7, 7, 'neigh_op_top_6')
// (7, 8, 'lutff_6/out')
// (7, 8, 'sp12_h_r_4')
// (7, 8, 'sp4_r_v_b_45')
// (7, 9, 'local_g0_3')
// (7, 9, 'lutff_4/in_1')
// (7, 9, 'neigh_op_bot_6')
// (7, 9, 'sp4_r_v_b_32')
// (7, 10, 'sp4_r_v_b_21')
// (7, 11, 'sp4_r_v_b_8')
// (8, 7, 'neigh_op_tnl_6')
// (8, 7, 'sp4_v_t_45')
// (8, 8, 'neigh_op_lft_6')
// (8, 8, 'sp12_h_r_7')
// (8, 8, 'sp4_v_b_45')
// (8, 9, 'neigh_op_bnl_6')
// (8, 9, 'sp4_v_b_32')
// (8, 10, 'sp4_v_b_21')
// (8, 11, 'sp4_v_b_8')
// (9, 8, 'sp12_h_r_8')
// (10, 8, 'sp12_h_r_11')
// (11, 8, 'local_g1_4')
// (11, 8, 'lutff_1/in_0')
// (11, 8, 'sp12_h_r_12')
// (12, 8, 'sp12_h_r_15')
// (13, 8, 'span12_horz_15')

reg n256 = 0;
// (5, 8, 'sp4_h_r_6')
// (6, 8, 'local_g0_3')
// (6, 8, 'lutff_6/in_1')
// (6, 8, 'sp4_h_r_19')
// (7, 8, 'sp4_h_r_30')
// (8, 8, 'sp4_h_r_43')
// (9, 8, 'sp4_h_l_43')
// (9, 8, 'sp4_h_r_10')
// (10, 7, 'neigh_op_tnr_1')
// (10, 8, 'neigh_op_rgt_1')
// (10, 8, 'sp4_h_r_23')
// (10, 9, 'neigh_op_bnr_1')
// (11, 7, 'neigh_op_top_1')
// (11, 8, 'lutff_1/out')
// (11, 8, 'sp4_h_r_34')
// (11, 9, 'neigh_op_bot_1')
// (12, 7, 'neigh_op_tnl_1')
// (12, 8, 'neigh_op_lft_1')
// (12, 8, 'sp4_h_r_47')
// (12, 9, 'neigh_op_bnl_1')
// (13, 8, 'span4_horz_47')

reg n257 = 0;
// (5, 9, 'neigh_op_tnr_0')
// (5, 10, 'neigh_op_rgt_0')
// (5, 11, 'neigh_op_bnr_0')
// (6, 7, 'sp4_r_v_b_36')
// (6, 8, 'sp4_r_v_b_25')
// (6, 9, 'neigh_op_top_0')
// (6, 9, 'sp4_r_v_b_12')
// (6, 10, 'lutff_0/out')
// (6, 10, 'sp4_r_v_b_1')
// (6, 11, 'local_g1_0')
// (6, 11, 'lutff_7/in_0')
// (6, 11, 'neigh_op_bot_0')
// (7, 6, 'sp4_h_r_1')
// (7, 6, 'sp4_v_t_36')
// (7, 7, 'sp4_v_b_36')
// (7, 8, 'sp4_v_b_25')
// (7, 9, 'neigh_op_tnl_0')
// (7, 9, 'sp4_v_b_12')
// (7, 10, 'neigh_op_lft_0')
// (7, 10, 'sp4_v_b_1')
// (7, 11, 'neigh_op_bnl_0')
// (8, 6, 'sp4_h_r_12')
// (9, 6, 'sp4_h_r_25')
// (10, 6, 'sp4_h_r_36')
// (10, 7, 'sp4_r_v_b_43')
// (10, 8, 'sp4_r_v_b_30')
// (10, 9, 'sp4_r_v_b_19')
// (10, 10, 'sp4_r_v_b_6')
// (11, 6, 'sp4_h_l_36')
// (11, 6, 'sp4_v_t_43')
// (11, 7, 'sp4_v_b_43')
// (11, 8, 'sp4_v_b_30')
// (11, 9, 'local_g0_3')
// (11, 9, 'lutff_0/in_3')
// (11, 9, 'lutff_3/in_0')
// (11, 9, 'sp4_v_b_19')
// (11, 10, 'sp4_v_b_6')

reg n258 = 0;
// (5, 9, 'neigh_op_tnr_1')
// (5, 10, 'neigh_op_rgt_1')
// (5, 11, 'neigh_op_bnr_1')
// (6, 9, 'neigh_op_top_1')
// (6, 10, 'local_g1_1')
// (6, 10, 'lutff_1/out')
// (6, 10, 'lutff_6/in_0')
// (6, 11, 'neigh_op_bot_1')
// (7, 9, 'neigh_op_tnl_1')
// (7, 10, 'neigh_op_lft_1')
// (7, 11, 'neigh_op_bnl_1')

reg n259 = 0;
// (5, 9, 'neigh_op_tnr_3')
// (5, 10, 'neigh_op_rgt_3')
// (5, 11, 'neigh_op_bnr_3')
// (6, 9, 'neigh_op_top_3')
// (6, 10, 'local_g1_3')
// (6, 10, 'lutff_3/out')
// (6, 10, 'lutff_5/in_3')
// (6, 11, 'neigh_op_bot_3')
// (7, 9, 'neigh_op_tnl_3')
// (7, 10, 'neigh_op_lft_3')
// (7, 11, 'neigh_op_bnl_3')

reg n260 = 0;
// (5, 9, 'neigh_op_tnr_4')
// (5, 10, 'neigh_op_rgt_4')
// (5, 11, 'neigh_op_bnr_4')
// (6, 9, 'neigh_op_top_4')
// (6, 10, 'local_g1_4')
// (6, 10, 'lutff_3/in_0')
// (6, 10, 'lutff_4/out')
// (6, 11, 'neigh_op_bot_4')
// (7, 9, 'neigh_op_tnl_4')
// (7, 10, 'neigh_op_lft_4')
// (7, 11, 'neigh_op_bnl_4')

reg n261 = 0;
// (5, 9, 'neigh_op_tnr_5')
// (5, 10, 'neigh_op_rgt_5')
// (5, 11, 'neigh_op_bnr_5')
// (6, 9, 'neigh_op_top_5')
// (6, 10, 'local_g0_5')
// (6, 10, 'lutff_1/in_0')
// (6, 10, 'lutff_5/out')
// (6, 11, 'neigh_op_bot_5')
// (7, 9, 'neigh_op_tnl_5')
// (7, 10, 'neigh_op_lft_5')
// (7, 11, 'neigh_op_bnl_5')

reg n262 = 0;
// (5, 9, 'neigh_op_tnr_6')
// (5, 10, 'neigh_op_rgt_6')
// (5, 11, 'neigh_op_bnr_6')
// (6, 9, 'neigh_op_top_6')
// (6, 10, 'local_g1_6')
// (6, 10, 'lutff_6/out')
// (6, 10, 'lutff_7/in_0')
// (6, 11, 'neigh_op_bot_6')
// (7, 9, 'neigh_op_tnl_6')
// (7, 10, 'neigh_op_lft_6')
// (7, 11, 'neigh_op_bnl_6')

reg n263 = 0;
// (5, 9, 'neigh_op_tnr_7')
// (5, 10, 'local_g3_7')
// (5, 10, 'lutff_5/in_3')
// (5, 10, 'neigh_op_rgt_7')
// (5, 11, 'local_g0_7')
// (5, 11, 'lutff_6/in_3')
// (5, 11, 'neigh_op_bnr_7')
// (6, 9, 'neigh_op_top_7')
// (6, 10, 'local_g2_7')
// (6, 10, 'lutff_5/in_2')
// (6, 10, 'lutff_7/out')
// (6, 11, 'neigh_op_bot_7')
// (7, 9, 'neigh_op_tnl_7')
// (7, 10, 'neigh_op_lft_7')
// (7, 11, 'neigh_op_bnl_7')

wire n264;
// (5, 9, 'sp4_h_r_2')
// (6, 8, 'neigh_op_tnr_5')
// (6, 9, 'neigh_op_rgt_5')
// (6, 9, 'sp4_h_r_15')
// (6, 10, 'neigh_op_bnr_5')
// (7, 8, 'neigh_op_top_5')
// (7, 9, 'lutff_5/out')
// (7, 9, 'sp4_h_r_26')
// (7, 10, 'local_g0_5')
// (7, 10, 'local_g1_5')
// (7, 10, 'lutff_4/in_1')
// (7, 10, 'lutff_5/in_3')
// (7, 10, 'neigh_op_bot_5')
// (8, 8, 'neigh_op_tnl_5')
// (8, 9, 'neigh_op_lft_5')
// (8, 9, 'sp4_h_r_39')
// (8, 10, 'neigh_op_bnl_5')
// (8, 10, 'sp4_r_v_b_42')
// (8, 11, 'sp4_r_v_b_31')
// (8, 12, 'sp4_r_v_b_18')
// (8, 13, 'sp4_r_v_b_7')
// (9, 9, 'sp4_h_l_39')
// (9, 9, 'sp4_v_t_42')
// (9, 10, 'local_g2_2')
// (9, 10, 'local_g3_2')
// (9, 10, 'lutff_1/in_1')
// (9, 10, 'lutff_3/in_2')
// (9, 10, 'lutff_4/in_1')
// (9, 10, 'lutff_5/in_3')
// (9, 10, 'lutff_6/in_3')
// (9, 10, 'lutff_7/in_3')
// (9, 10, 'sp4_v_b_42')
// (9, 11, 'sp4_v_b_31')
// (9, 12, 'sp4_v_b_18')
// (9, 13, 'sp4_v_b_7')

wire n265;
// (5, 9, 'sp4_r_v_b_36')
// (5, 10, 'neigh_op_tnr_6')
// (5, 10, 'sp4_r_v_b_25')
// (5, 11, 'neigh_op_rgt_6')
// (5, 11, 'sp4_r_v_b_12')
// (5, 12, 'neigh_op_bnr_6')
// (5, 12, 'sp4_r_v_b_1')
// (6, 8, 'sp4_v_t_36')
// (6, 9, 'sp4_v_b_36')
// (6, 10, 'neigh_op_top_6')
// (6, 10, 'sp4_v_b_25')
// (6, 11, 'lutff_6/out')
// (6, 11, 'sp4_v_b_12')
// (6, 12, 'local_g1_1')
// (6, 12, 'local_g1_6')
// (6, 12, 'lutff_0/in_0')
// (6, 12, 'lutff_1/in_2')
// (6, 12, 'neigh_op_bot_6')
// (6, 12, 'sp4_v_b_1')
// (7, 10, 'neigh_op_tnl_6')
// (7, 11, 'neigh_op_lft_6')
// (7, 12, 'neigh_op_bnl_6')

wire n266;
// (5, 10, 'neigh_op_tnr_1')
// (5, 11, 'neigh_op_rgt_1')
// (5, 12, 'neigh_op_bnr_1')
// (6, 10, 'neigh_op_top_1')
// (6, 11, 'local_g0_1')
// (6, 11, 'local_g3_1')
// (6, 11, 'lutff_1/out')
// (6, 11, 'lutff_2/in_1')
// (6, 11, 'lutff_4/in_2')
// (6, 12, 'neigh_op_bot_1')
// (7, 10, 'neigh_op_tnl_1')
// (7, 11, 'neigh_op_lft_1')
// (7, 12, 'neigh_op_bnl_1')

wire n267;
// (5, 10, 'neigh_op_tnr_2')
// (5, 11, 'neigh_op_rgt_2')
// (5, 12, 'neigh_op_bnr_2')
// (6, 1, 'sp12_v_t_23')
// (6, 2, 'sp12_v_b_23')
// (6, 3, 'sp12_v_b_20')
// (6, 4, 'sp12_v_b_19')
// (6, 5, 'sp12_v_b_16')
// (6, 6, 'sp12_v_b_15')
// (6, 7, 'sp12_v_b_12')
// (6, 8, 'sp12_v_b_11')
// (6, 9, 'sp12_v_b_8')
// (6, 10, 'neigh_op_top_2')
// (6, 10, 'sp12_v_b_7')
// (6, 11, 'lutff_2/out')
// (6, 11, 'sp12_v_b_4')
// (6, 12, 'local_g2_3')
// (6, 12, 'lutff_2/in_3')
// (6, 12, 'lutff_5/in_2')
// (6, 12, 'lutff_6/in_1')
// (6, 12, 'neigh_op_bot_2')
// (6, 12, 'sp12_v_b_3')
// (6, 13, 'sp12_v_b_0')
// (7, 10, 'neigh_op_tnl_2')
// (7, 11, 'neigh_op_lft_2')
// (7, 12, 'neigh_op_bnl_2')

wire n268;
// (5, 10, 'neigh_op_tnr_3')
// (5, 11, 'neigh_op_rgt_3')
// (5, 12, 'neigh_op_bnr_3')
// (6, 10, 'neigh_op_top_3')
// (6, 11, 'lutff_3/out')
// (6, 11, 'sp4_r_v_b_39')
// (6, 12, 'local_g1_2')
// (6, 12, 'local_g1_3')
// (6, 12, 'lutff_0/in_3')
// (6, 12, 'lutff_1/in_3')
// (6, 12, 'neigh_op_bot_3')
// (6, 12, 'sp4_r_v_b_26')
// (6, 13, 'sp4_r_v_b_15')
// (6, 14, 'sp4_r_v_b_2')
// (7, 10, 'neigh_op_tnl_3')
// (7, 10, 'sp4_v_t_39')
// (7, 11, 'neigh_op_lft_3')
// (7, 11, 'sp4_v_b_39')
// (7, 12, 'neigh_op_bnl_3')
// (7, 12, 'sp4_v_b_26')
// (7, 13, 'sp4_v_b_15')
// (7, 14, 'sp4_v_b_2')

wire n269;
// (5, 10, 'neigh_op_tnr_4')
// (5, 11, 'neigh_op_rgt_4')
// (5, 11, 'sp4_r_v_b_40')
// (5, 12, 'neigh_op_bnr_4')
// (5, 12, 'sp4_r_v_b_29')
// (5, 13, 'sp4_r_v_b_16')
// (5, 14, 'sp4_r_v_b_5')
// (6, 3, 'sp12_v_t_23')
// (6, 4, 'sp12_v_b_23')
// (6, 5, 'sp12_v_b_20')
// (6, 6, 'sp12_v_b_19')
// (6, 7, 'sp12_v_b_16')
// (6, 8, 'sp12_v_b_15')
// (6, 9, 'sp12_v_b_12')
// (6, 10, 'neigh_op_top_4')
// (6, 10, 'sp12_v_b_11')
// (6, 10, 'sp4_v_t_40')
// (6, 11, 'lutff_4/out')
// (6, 11, 'sp12_v_b_8')
// (6, 11, 'sp4_v_b_40')
// (6, 12, 'local_g3_5')
// (6, 12, 'lutff_4/in_2')
// (6, 12, 'neigh_op_bot_4')
// (6, 12, 'sp12_v_b_7')
// (6, 12, 'sp4_v_b_29')
// (6, 13, 'local_g1_0')
// (6, 13, 'local_g2_4')
// (6, 13, 'lutff_4/in_2')
// (6, 13, 'lutff_5/in_3')
// (6, 13, 'lutff_6/in_1')
// (6, 13, 'sp12_v_b_4')
// (6, 13, 'sp4_v_b_16')
// (6, 14, 'sp12_v_b_3')
// (6, 14, 'sp4_v_b_5')
// (6, 15, 'sp12_v_b_0')
// (7, 10, 'neigh_op_tnl_4')
// (7, 11, 'neigh_op_lft_4')
// (7, 12, 'neigh_op_bnl_4')

reg n270 = 0;
// (5, 10, 'neigh_op_tnr_7')
// (5, 11, 'neigh_op_rgt_7')
// (5, 12, 'neigh_op_bnr_7')
// (6, 10, 'neigh_op_top_7')
// (6, 11, 'local_g3_7')
// (6, 11, 'lutff_3/in_3')
// (6, 11, 'lutff_7/out')
// (6, 12, 'neigh_op_bot_7')
// (7, 10, 'neigh_op_tnl_7')
// (7, 11, 'neigh_op_lft_7')
// (7, 12, 'neigh_op_bnl_7')

wire n271;
// (5, 11, 'neigh_op_tnr_0')
// (5, 12, 'neigh_op_rgt_0')
// (5, 13, 'neigh_op_bnr_0')
// (6, 11, 'neigh_op_top_0')
// (6, 11, 'sp4_r_v_b_44')
// (6, 12, 'local_g0_2')
// (6, 12, 'local_g1_0')
// (6, 12, 'lutff_0/out')
// (6, 12, 'lutff_4/in_3')
// (6, 12, 'lutff_5/in_3')
// (6, 12, 'sp4_r_v_b_33')
// (6, 13, 'neigh_op_bot_0')
// (6, 13, 'sp4_r_v_b_20')
// (6, 14, 'sp4_r_v_b_9')
// (7, 10, 'sp4_v_t_44')
// (7, 11, 'neigh_op_tnl_0')
// (7, 11, 'sp4_v_b_44')
// (7, 12, 'neigh_op_lft_0')
// (7, 12, 'sp4_v_b_33')
// (7, 13, 'neigh_op_bnl_0')
// (7, 13, 'sp4_v_b_20')
// (7, 14, 'sp4_v_b_9')

wire n272;
// (5, 11, 'neigh_op_tnr_1')
// (5, 11, 'sp4_r_v_b_47')
// (5, 12, 'neigh_op_rgt_1')
// (5, 12, 'sp4_r_v_b_34')
// (5, 13, 'neigh_op_bnr_1')
// (5, 13, 'sp4_r_v_b_23')
// (5, 14, 'sp4_r_v_b_10')
// (6, 10, 'sp4_v_t_47')
// (6, 11, 'neigh_op_top_1')
// (6, 11, 'sp4_v_b_47')
// (6, 12, 'local_g3_2')
// (6, 12, 'lutff_1/out')
// (6, 12, 'lutff_6/in_3')
// (6, 12, 'sp4_v_b_34')
// (6, 13, 'neigh_op_bot_1')
// (6, 13, 'sp4_v_b_23')
// (6, 14, 'sp4_v_b_10')
// (7, 11, 'neigh_op_tnl_1')
// (7, 12, 'neigh_op_lft_1')
// (7, 13, 'neigh_op_bnl_1')

wire n273;
// (5, 11, 'neigh_op_tnr_2')
// (5, 12, 'neigh_op_rgt_2')
// (5, 12, 'sp4_r_v_b_36')
// (5, 13, 'neigh_op_bnr_2')
// (5, 13, 'sp4_r_v_b_25')
// (5, 14, 'sp4_r_v_b_12')
// (5, 15, 'sp4_r_v_b_1')
// (6, 2, 'sp12_v_t_23')
// (6, 3, 'sp12_v_b_23')
// (6, 4, 'sp12_v_b_20')
// (6, 5, 'sp12_v_b_19')
// (6, 6, 'sp12_v_b_16')
// (6, 7, 'sp12_v_b_15')
// (6, 8, 'sp12_v_b_12')
// (6, 9, 'sp12_v_b_11')
// (6, 10, 'sp12_v_b_8')
// (6, 11, 'neigh_op_top_2')
// (6, 11, 'sp12_v_b_7')
// (6, 11, 'sp4_v_t_36')
// (6, 12, 'lutff_2/out')
// (6, 12, 'sp12_v_b_4')
// (6, 12, 'sp4_v_b_36')
// (6, 13, 'neigh_op_bot_2')
// (6, 13, 'sp12_v_b_3')
// (6, 13, 'sp4_v_b_25')
// (6, 14, 'local_g1_4')
// (6, 14, 'local_g2_0')
// (6, 14, 'lutff_0/in_1')
// (6, 14, 'lutff_1/in_3')
// (6, 14, 'lutff_2/in_3')
// (6, 14, 'sp12_v_b_0')
// (6, 14, 'sp4_v_b_12')
// (6, 15, 'sp4_v_b_1')
// (7, 11, 'neigh_op_tnl_2')
// (7, 12, 'neigh_op_lft_2')
// (7, 13, 'neigh_op_bnl_2')

wire n274;
// (5, 11, 'neigh_op_tnr_7')
// (5, 11, 'sp4_r_v_b_43')
// (5, 12, 'neigh_op_rgt_7')
// (5, 12, 'sp4_r_v_b_30')
// (5, 12, 'sp4_r_v_b_46')
// (5, 13, 'neigh_op_bnr_7')
// (5, 13, 'sp4_r_v_b_19')
// (5, 13, 'sp4_r_v_b_35')
// (5, 14, 'sp4_r_v_b_22')
// (5, 14, 'sp4_r_v_b_6')
// (5, 15, 'sp4_r_v_b_11')
// (6, 10, 'sp4_v_t_43')
// (6, 11, 'neigh_op_top_7')
// (6, 11, 'sp4_v_b_43')
// (6, 11, 'sp4_v_t_46')
// (6, 12, 'lutff_7/out')
// (6, 12, 'sp4_v_b_30')
// (6, 12, 'sp4_v_b_46')
// (6, 13, 'neigh_op_bot_7')
// (6, 13, 'sp4_v_b_19')
// (6, 13, 'sp4_v_b_35')
// (6, 14, 'local_g0_6')
// (6, 14, 'lutff_5/in_3')
// (6, 14, 'sp4_h_r_6')
// (6, 14, 'sp4_v_b_22')
// (6, 14, 'sp4_v_b_6')
// (6, 15, 'local_g0_3')
// (6, 15, 'local_g1_3')
// (6, 15, 'lutff_0/in_2')
// (6, 15, 'lutff_7/in_2')
// (6, 15, 'sp4_h_r_5')
// (6, 15, 'sp4_v_b_11')
// (7, 11, 'neigh_op_tnl_7')
// (7, 12, 'neigh_op_lft_7')
// (7, 13, 'neigh_op_bnl_7')
// (7, 14, 'local_g1_3')
// (7, 14, 'lutff_0/in_2')
// (7, 14, 'sp4_h_r_19')
// (7, 15, 'local_g1_0')
// (7, 15, 'lutff_2/in_3')
// (7, 15, 'sp4_h_r_16')
// (8, 14, 'sp4_h_r_30')
// (8, 15, 'sp4_h_r_29')
// (9, 14, 'sp4_h_r_43')
// (9, 15, 'sp4_h_r_40')
// (10, 14, 'sp4_h_l_43')
// (10, 15, 'sp4_h_l_40')

wire n275;
// (5, 11, 'sp4_h_r_7')
// (6, 11, 'sp4_h_r_18')
// (7, 10, 'neigh_op_tnr_5')
// (7, 11, 'neigh_op_rgt_5')
// (7, 11, 'sp4_h_r_31')
// (7, 12, 'neigh_op_bnr_5')
// (8, 10, 'neigh_op_top_5')
// (8, 11, 'local_g0_5')
// (8, 11, 'local_g2_2')
// (8, 11, 'lutff_1/in_3')
// (8, 11, 'lutff_2/in_3')
// (8, 11, 'lutff_5/out')
// (8, 11, 'sp4_h_r_42')
// (8, 12, 'neigh_op_bot_5')
// (9, 10, 'neigh_op_tnl_5')
// (9, 11, 'neigh_op_lft_5')
// (9, 11, 'sp4_h_l_42')
// (9, 12, 'neigh_op_bnl_5')

wire n276;
// (5, 12, 'neigh_op_tnr_0')
// (5, 13, 'neigh_op_rgt_0')
// (5, 14, 'neigh_op_bnr_0')
// (6, 10, 'sp4_r_v_b_36')
// (6, 11, 'sp4_r_v_b_25')
// (6, 12, 'neigh_op_top_0')
// (6, 12, 'sp4_r_v_b_12')
// (6, 13, 'local_g0_0')
// (6, 13, 'lutff_0/out')
// (6, 13, 'lutff_4/in_0')
// (6, 13, 'lutff_6/in_0')
// (6, 13, 'sp4_r_v_b_1')
// (6, 14, 'neigh_op_bot_0')
// (7, 9, 'sp4_v_t_36')
// (7, 10, 'sp4_v_b_36')
// (7, 11, 'sp4_v_b_25')
// (7, 12, 'neigh_op_tnl_0')
// (7, 12, 'sp4_v_b_12')
// (7, 13, 'local_g1_1')
// (7, 13, 'lutff_0/in_2')
// (7, 13, 'lutff_3/in_3')
// (7, 13, 'neigh_op_lft_0')
// (7, 13, 'sp4_v_b_1')
// (7, 14, 'neigh_op_bnl_0')

wire n277;
// (5, 12, 'neigh_op_tnr_2')
// (5, 13, 'neigh_op_rgt_2')
// (5, 14, 'neigh_op_bnr_2')
// (6, 12, 'neigh_op_top_2')
// (6, 13, 'local_g0_2')
// (6, 13, 'local_g1_2')
// (6, 13, 'lutff_2/out')
// (6, 13, 'lutff_4/in_3')
// (6, 13, 'lutff_6/in_2')
// (6, 14, 'local_g1_2')
// (6, 14, 'lutff_2/in_1')
// (6, 14, 'neigh_op_bot_2')
// (7, 12, 'neigh_op_tnl_2')
// (7, 13, 'local_g0_2')
// (7, 13, 'local_g1_2')
// (7, 13, 'lutff_1/in_1')
// (7, 13, 'lutff_4/in_3')
// (7, 13, 'neigh_op_lft_2')
// (7, 14, 'neigh_op_bnl_2')

wire n278;
// (5, 12, 'neigh_op_tnr_3')
// (5, 13, 'neigh_op_rgt_3')
// (5, 13, 'sp4_h_r_11')
// (5, 14, 'neigh_op_bnr_3')
// (6, 12, 'neigh_op_top_3')
// (6, 13, 'lutff_3/out')
// (6, 13, 'sp4_h_r_22')
// (6, 14, 'local_g0_3')
// (6, 14, 'local_g1_3')
// (6, 14, 'lutff_0/in_3')
// (6, 14, 'lutff_1/in_2')
// (6, 14, 'lutff_2/in_2')
// (6, 14, 'lutff_6/in_3')
// (6, 14, 'neigh_op_bot_3')
// (7, 12, 'neigh_op_tnl_3')
// (7, 13, 'neigh_op_lft_3')
// (7, 13, 'sp4_h_r_35')
// (7, 14, 'neigh_op_bnl_3')
// (8, 13, 'sp4_h_r_46')
// (8, 14, 'local_g3_1')
// (8, 14, 'lutff_3/in_1')
// (8, 14, 'lutff_5/in_1')
// (8, 14, 'lutff_6/in_2')
// (8, 14, 'sp4_r_v_b_41')
// (8, 15, 'sp4_r_v_b_28')
// (8, 16, 'sp4_r_v_b_17')
// (9, 13, 'sp4_h_l_46')
// (9, 13, 'sp4_v_t_41')
// (9, 14, 'sp4_v_b_41')
// (9, 15, 'sp4_v_b_28')
// (9, 16, 'sp4_v_b_17')
// (9, 17, 'span4_vert_4')

wire n279;
// (5, 12, 'neigh_op_tnr_4')
// (5, 13, 'neigh_op_rgt_4')
// (5, 14, 'neigh_op_bnr_4')
// (6, 12, 'neigh_op_top_4')
// (6, 13, 'lutff_4/out')
// (6, 14, 'local_g0_4')
// (6, 14, 'lutff_7/in_3')
// (6, 14, 'neigh_op_bot_4')
// (7, 12, 'neigh_op_tnl_4')
// (7, 13, 'neigh_op_lft_4')
// (7, 14, 'neigh_op_bnl_4')

wire n280;
// (5, 12, 'neigh_op_tnr_5')
// (5, 13, 'neigh_op_rgt_5')
// (5, 14, 'neigh_op_bnr_5')
// (6, 10, 'sp4_r_v_b_46')
// (6, 11, 'sp4_r_v_b_35')
// (6, 12, 'neigh_op_top_5')
// (6, 12, 'sp4_r_v_b_22')
// (6, 13, 'lutff_5/out')
// (6, 13, 'sp4_h_r_10')
// (6, 13, 'sp4_r_v_b_11')
// (6, 14, 'neigh_op_bot_5')
// (7, 9, 'sp4_v_t_46')
// (7, 10, 'sp4_v_b_46')
// (7, 11, 'sp4_v_b_35')
// (7, 12, 'neigh_op_tnl_5')
// (7, 12, 'sp4_v_b_22')
// (7, 13, 'local_g0_5')
// (7, 13, 'local_g1_3')
// (7, 13, 'lutff_0/in_1')
// (7, 13, 'lutff_2/in_2')
// (7, 13, 'lutff_3/in_1')
// (7, 13, 'neigh_op_lft_5')
// (7, 13, 'sp4_h_r_23')
// (7, 13, 'sp4_v_b_11')
// (7, 14, 'neigh_op_bnl_5')
// (8, 13, 'local_g3_2')
// (8, 13, 'lutff_5/in_2')
// (8, 13, 'sp4_h_r_34')
// (9, 13, 'sp4_h_r_47')
// (10, 13, 'sp4_h_l_47')

wire n281;
// (5, 12, 'neigh_op_tnr_6')
// (5, 12, 'sp4_r_v_b_41')
// (5, 13, 'neigh_op_rgt_6')
// (5, 13, 'sp4_r_v_b_28')
// (5, 14, 'neigh_op_bnr_6')
// (5, 14, 'sp4_r_v_b_17')
// (5, 15, 'sp4_r_v_b_4')
// (6, 11, 'sp4_v_t_41')
// (6, 12, 'neigh_op_top_6')
// (6, 12, 'sp4_v_b_41')
// (6, 13, 'lutff_6/out')
// (6, 13, 'sp4_v_b_28')
// (6, 14, 'neigh_op_bot_6')
// (6, 14, 'sp4_v_b_17')
// (6, 15, 'local_g0_4')
// (6, 15, 'lutff_3/in_3')
// (6, 15, 'sp4_v_b_4')
// (7, 12, 'neigh_op_tnl_6')
// (7, 13, 'neigh_op_lft_6')
// (7, 14, 'neigh_op_bnl_6')

wire n282;
// (5, 12, 'neigh_op_tnr_7')
// (5, 13, 'neigh_op_rgt_7')
// (5, 14, 'neigh_op_bnr_7')
// (6, 12, 'neigh_op_top_7')
// (6, 13, 'lutff_7/out')
// (6, 14, 'local_g0_7')
// (6, 14, 'lutff_4/in_3')
// (6, 14, 'lutff_5/in_2')
// (6, 14, 'neigh_op_bot_7')
// (7, 12, 'neigh_op_tnl_7')
// (7, 13, 'neigh_op_lft_7')
// (7, 14, 'local_g2_7')
// (7, 14, 'lutff_5/in_2')
// (7, 14, 'neigh_op_bnl_7')

wire n283;
// (5, 12, 'sp4_h_r_10')
// (6, 11, 'neigh_op_tnr_1')
// (6, 12, 'local_g0_7')
// (6, 12, 'lutff_3/in_2')
// (6, 12, 'neigh_op_rgt_1')
// (6, 12, 'sp4_h_r_23')
// (6, 13, 'neigh_op_bnr_1')
// (7, 11, 'neigh_op_top_1')
// (7, 12, 'lutff_1/out')
// (7, 12, 'sp4_h_r_34')
// (7, 13, 'neigh_op_bot_1')
// (8, 11, 'neigh_op_tnl_1')
// (8, 12, 'neigh_op_lft_1')
// (8, 12, 'sp4_h_r_47')
// (8, 13, 'neigh_op_bnl_1')
// (9, 12, 'sp4_h_l_47')

wire n284;
// (5, 13, 'neigh_op_tnr_0')
// (5, 14, 'neigh_op_rgt_0')
// (5, 15, 'neigh_op_bnr_0')
// (6, 10, 'sp12_v_t_23')
// (6, 11, 'sp12_v_b_23')
// (6, 12, 'sp12_v_b_20')
// (6, 13, 'neigh_op_top_0')
// (6, 13, 'sp12_v_b_19')
// (6, 14, 'lutff_0/out')
// (6, 14, 'sp12_v_b_16')
// (6, 15, 'local_g3_7')
// (6, 15, 'lutff_7/in_3')
// (6, 15, 'neigh_op_bot_0')
// (6, 15, 'sp12_v_b_15')
// (6, 16, 'sp12_v_b_12')
// (6, 17, 'span12_vert_11')
// (7, 13, 'neigh_op_tnl_0')
// (7, 14, 'neigh_op_lft_0')
// (7, 15, 'neigh_op_bnl_0')

wire n285;
// (5, 13, 'neigh_op_tnr_1')
// (5, 14, 'neigh_op_rgt_1')
// (5, 15, 'neigh_op_bnr_1')
// (6, 11, 'sp4_r_v_b_38')
// (6, 12, 'sp4_r_v_b_27')
// (6, 13, 'neigh_op_top_1')
// (6, 13, 'sp4_r_v_b_14')
// (6, 14, 'lutff_1/out')
// (6, 14, 'sp4_r_v_b_3')
// (6, 15, 'local_g0_1')
// (6, 15, 'local_g1_1')
// (6, 15, 'lutff_0/in_1')
// (6, 15, 'lutff_7/in_1')
// (6, 15, 'neigh_op_bot_1')
// (7, 10, 'sp4_v_t_38')
// (7, 11, 'sp4_v_b_38')
// (7, 12, 'sp4_v_b_27')
// (7, 13, 'neigh_op_tnl_1')
// (7, 13, 'sp4_v_b_14')
// (7, 14, 'local_g0_3')
// (7, 14, 'lutff_3/in_0')
// (7, 14, 'neigh_op_lft_1')
// (7, 14, 'sp4_v_b_3')
// (7, 15, 'local_g3_1')
// (7, 15, 'lutff_2/in_2')
// (7, 15, 'neigh_op_bnl_1')

wire n286;
// (5, 13, 'neigh_op_tnr_4')
// (5, 14, 'neigh_op_rgt_4')
// (5, 15, 'neigh_op_bnr_4')
// (6, 13, 'neigh_op_top_4')
// (6, 14, 'lutff_4/out')
// (6, 15, 'local_g1_4')
// (6, 15, 'lutff_0/in_3')
// (6, 15, 'lutff_7/in_0')
// (6, 15, 'neigh_op_bot_4')
// (7, 13, 'neigh_op_tnl_4')
// (7, 14, 'neigh_op_lft_4')
// (7, 15, 'local_g2_4')
// (7, 15, 'lutff_1/in_3')
// (7, 15, 'neigh_op_bnl_4')

wire n287;
// (5, 13, 'neigh_op_tnr_5')
// (5, 14, 'neigh_op_rgt_5')
// (5, 15, 'neigh_op_bnr_5')
// (6, 13, 'neigh_op_top_5')
// (6, 14, 'lutff_5/out')
// (6, 15, 'local_g0_5')
// (6, 15, 'local_g1_5')
// (6, 15, 'lutff_1/in_1')
// (6, 15, 'lutff_2/in_1')
// (6, 15, 'neigh_op_bot_5')
// (7, 13, 'neigh_op_tnl_5')
// (7, 14, 'neigh_op_lft_5')
// (7, 15, 'neigh_op_bnl_5')

wire n288;
// (5, 13, 'neigh_op_tnr_6')
// (5, 14, 'neigh_op_rgt_6')
// (5, 15, 'neigh_op_bnr_6')
// (6, 13, 'neigh_op_top_6')
// (6, 14, 'local_g1_6')
// (6, 14, 'lutff_6/out')
// (6, 14, 'lutff_7/in_2')
// (6, 15, 'local_g0_6')
// (6, 15, 'local_g1_6')
// (6, 15, 'lutff_1/in_3')
// (6, 15, 'lutff_2/in_3')
// (6, 15, 'lutff_3/in_2')
// (6, 15, 'neigh_op_bot_6')
// (7, 13, 'neigh_op_tnl_6')
// (7, 14, 'neigh_op_lft_6')
// (7, 15, 'neigh_op_bnl_6')

wire n289;
// (5, 14, 'neigh_op_tnr_0')
// (5, 15, 'neigh_op_rgt_0')
// (5, 16, 'neigh_op_bnr_0')
// (6, 14, 'neigh_op_top_0')
// (6, 15, 'local_g0_0')
// (6, 15, 'local_g1_0')
// (6, 15, 'lutff_0/out')
// (6, 15, 'lutff_1/in_2')
// (6, 15, 'lutff_2/in_2')
// (6, 16, 'neigh_op_bot_0')
// (7, 14, 'neigh_op_tnl_0')
// (7, 15, 'neigh_op_lft_0')
// (7, 16, 'neigh_op_bnl_0')

wire n290;
// (5, 14, 'neigh_op_tnr_2')
// (5, 15, 'neigh_op_rgt_2')
// (5, 16, 'neigh_op_bnr_2')
// (6, 14, 'neigh_op_top_2')
// (6, 15, 'lutff_2/out')
// (6, 16, 'neigh_op_bot_2')
// (7, 14, 'neigh_op_tnl_2')
// (7, 15, 'local_g1_2')
// (7, 15, 'lutff_1/in_0')
// (7, 15, 'lutff_7/in_0')
// (7, 15, 'neigh_op_lft_2')
// (7, 16, 'neigh_op_bnl_2')

wire n291;
// (5, 14, 'neigh_op_tnr_3')
// (5, 15, 'neigh_op_rgt_3')
// (5, 15, 'sp4_h_r_11')
// (5, 16, 'neigh_op_bnr_3')
// (6, 14, 'neigh_op_top_3')
// (6, 15, 'lutff_3/out')
// (6, 15, 'sp4_h_r_22')
// (6, 16, 'neigh_op_bot_3')
// (7, 14, 'neigh_op_tnl_3')
// (7, 15, 'local_g2_3')
// (7, 15, 'lutff_4/in_3')
// (7, 15, 'lutff_6/in_3')
// (7, 15, 'neigh_op_lft_3')
// (7, 15, 'sp4_h_r_35')
// (7, 16, 'neigh_op_bnl_3')
// (8, 15, 'sp4_h_r_46')
// (9, 15, 'sp4_h_l_46')

wire n292;
// (5, 14, 'neigh_op_tnr_7')
// (5, 15, 'neigh_op_rgt_7')
// (5, 16, 'neigh_op_bnr_7')
// (6, 14, 'neigh_op_top_7')
// (6, 15, 'lutff_7/out')
// (6, 16, 'neigh_op_bot_7')
// (7, 14, 'neigh_op_tnl_7')
// (7, 15, 'local_g0_7')
// (7, 15, 'local_g1_7')
// (7, 15, 'lutff_0/in_3')
// (7, 15, 'lutff_6/in_2')
// (7, 15, 'neigh_op_lft_7')
// (7, 16, 'neigh_op_bnl_7')

wire n293;
// (5, 14, 'sp4_h_r_11')
// (6, 14, 'sp4_h_r_22')
// (7, 13, 'local_g2_7')
// (7, 13, 'local_g3_7')
// (7, 13, 'lutff_5/in_2')
// (7, 13, 'lutff_7/in_1')
// (7, 13, 'neigh_op_tnr_7')
// (7, 14, 'local_g2_3')
// (7, 14, 'lutff_3/in_2')
// (7, 14, 'neigh_op_rgt_7')
// (7, 14, 'sp4_h_r_35')
// (7, 15, 'neigh_op_bnr_7')
// (8, 13, 'neigh_op_top_7')
// (8, 14, 'lutff_7/out')
// (8, 14, 'sp4_h_r_46')
// (8, 15, 'neigh_op_bot_7')
// (9, 13, 'neigh_op_tnl_7')
// (9, 14, 'neigh_op_lft_7')
// (9, 14, 'sp4_h_l_46')
// (9, 15, 'neigh_op_bnl_7')

reg n294 = 0;
// (6, 2, 'neigh_op_tnr_0')
// (6, 3, 'neigh_op_rgt_0')
// (6, 4, 'neigh_op_bnr_0')
// (7, 2, 'neigh_op_top_0')
// (7, 3, 'local_g1_0')
// (7, 3, 'lutff_0/out')
// (7, 3, 'lutff_1/in_0')
// (7, 4, 'neigh_op_bot_0')
// (8, 2, 'neigh_op_tnl_0')
// (8, 3, 'neigh_op_lft_0')
// (8, 4, 'neigh_op_bnl_0')

reg n295 = 0;
// (6, 2, 'neigh_op_tnr_1')
// (6, 3, 'neigh_op_rgt_1')
// (6, 4, 'neigh_op_bnr_1')
// (7, 2, 'neigh_op_top_1')
// (7, 3, 'lutff_1/out')
// (7, 4, 'local_g0_1')
// (7, 4, 'lutff_3/in_0')
// (7, 4, 'neigh_op_bot_1')
// (8, 2, 'neigh_op_tnl_1')
// (8, 3, 'neigh_op_lft_1')
// (8, 4, 'neigh_op_bnl_1')

reg n296 = 0;
// (6, 2, 'neigh_op_tnr_2')
// (6, 3, 'neigh_op_rgt_2')
// (6, 4, 'neigh_op_bnr_2')
// (7, 2, 'neigh_op_top_2')
// (7, 3, 'local_g0_2')
// (7, 3, 'lutff_2/out')
// (7, 3, 'lutff_4/in_0')
// (7, 4, 'neigh_op_bot_2')
// (8, 2, 'neigh_op_tnl_2')
// (8, 3, 'neigh_op_lft_2')
// (8, 4, 'neigh_op_bnl_2')

reg n297 = 0;
// (6, 2, 'neigh_op_tnr_3')
// (6, 3, 'neigh_op_rgt_3')
// (6, 4, 'neigh_op_bnr_3')
// (7, 2, 'neigh_op_top_3')
// (7, 3, 'local_g1_3')
// (7, 3, 'lutff_2/in_0')
// (7, 3, 'lutff_3/out')
// (7, 4, 'local_g0_3')
// (7, 4, 'local_g1_3')
// (7, 4, 'lutff_1/in_1')
// (7, 4, 'lutff_5/in_0')
// (7, 4, 'lutff_6/in_2')
// (7, 4, 'neigh_op_bot_3')
// (8, 2, 'neigh_op_tnl_3')
// (8, 3, 'neigh_op_lft_3')
// (8, 4, 'neigh_op_bnl_3')

reg n298 = 0;
// (6, 2, 'neigh_op_tnr_4')
// (6, 3, 'neigh_op_rgt_4')
// (6, 4, 'neigh_op_bnr_4')
// (7, 2, 'neigh_op_top_4')
// (7, 3, 'local_g0_4')
// (7, 3, 'lutff_4/out')
// (7, 3, 'lutff_6/in_0')
// (7, 4, 'neigh_op_bot_4')
// (8, 2, 'neigh_op_tnl_4')
// (8, 3, 'neigh_op_lft_4')
// (8, 4, 'neigh_op_bnl_4')

reg n299 = 0;
// (6, 2, 'neigh_op_tnr_6')
// (6, 3, 'neigh_op_rgt_6')
// (6, 4, 'neigh_op_bnr_6')
// (7, 2, 'neigh_op_top_6')
// (7, 3, 'local_g1_6')
// (7, 3, 'lutff_3/in_0')
// (7, 3, 'lutff_6/out')
// (7, 4, 'neigh_op_bot_6')
// (8, 2, 'neigh_op_tnl_6')
// (8, 3, 'neigh_op_lft_6')
// (8, 4, 'neigh_op_bnl_6')

wire n300;
// (6, 3, 'neigh_op_tnr_1')
// (6, 4, 'neigh_op_rgt_1')
// (6, 5, 'neigh_op_bnr_1')
// (7, 3, 'neigh_op_top_1')
// (7, 4, 'local_g2_1')
// (7, 4, 'lutff_0/in_3')
// (7, 4, 'lutff_1/out')
// (7, 5, 'neigh_op_bot_1')
// (8, 3, 'neigh_op_tnl_1')
// (8, 4, 'neigh_op_lft_1')
// (8, 5, 'neigh_op_bnl_1')

reg n301 = 0;
// (6, 3, 'neigh_op_tnr_2')
// (6, 4, 'neigh_op_rgt_2')
// (6, 5, 'neigh_op_bnr_2')
// (7, 3, 'neigh_op_top_2')
// (7, 4, 'local_g3_2')
// (7, 4, 'lutff_2/out')
// (7, 4, 'lutff_7/in_0')
// (7, 5, 'neigh_op_bot_2')
// (8, 3, 'neigh_op_tnl_2')
// (8, 4, 'neigh_op_lft_2')
// (8, 5, 'neigh_op_bnl_2')

reg n302 = 0;
// (6, 3, 'neigh_op_tnr_3')
// (6, 4, 'neigh_op_rgt_3')
// (6, 5, 'neigh_op_bnr_3')
// (7, 3, 'neigh_op_top_3')
// (7, 4, 'local_g2_3')
// (7, 4, 'local_g3_3')
// (7, 4, 'lutff_1/in_0')
// (7, 4, 'lutff_3/out')
// (7, 4, 'lutff_5/in_1')
// (7, 5, 'neigh_op_bot_3')
// (8, 3, 'neigh_op_tnl_3')
// (8, 4, 'neigh_op_lft_3')
// (8, 5, 'neigh_op_bnl_3')

reg n303 = 0;
// (6, 3, 'neigh_op_tnr_4')
// (6, 4, 'neigh_op_rgt_4')
// (6, 5, 'neigh_op_bnr_4')
// (7, 3, 'neigh_op_top_4')
// (7, 4, 'local_g0_4')
// (7, 4, 'lutff_2/in_0')
// (7, 4, 'lutff_4/out')
// (7, 5, 'neigh_op_bot_4')
// (8, 3, 'neigh_op_tnl_4')
// (8, 4, 'neigh_op_lft_4')
// (8, 5, 'neigh_op_bnl_4')

reg n304 = 0;
// (6, 3, 'neigh_op_tnr_5')
// (6, 4, 'neigh_op_rgt_5')
// (6, 5, 'neigh_op_bnr_5')
// (7, 3, 'neigh_op_top_5')
// (7, 4, 'local_g1_5')
// (7, 4, 'lutff_4/in_0')
// (7, 4, 'lutff_5/out')
// (7, 5, 'neigh_op_bot_5')
// (8, 3, 'neigh_op_tnl_5')
// (8, 4, 'neigh_op_lft_5')
// (8, 5, 'neigh_op_bnl_5')

reg n305 = 0;
// (6, 3, 'neigh_op_tnr_6')
// (6, 4, 'neigh_op_rgt_6')
// (6, 5, 'neigh_op_bnr_6')
// (7, 3, 'local_g0_6')
// (7, 3, 'lutff_0/in_0')
// (7, 3, 'neigh_op_top_6')
// (7, 4, 'lutff_6/out')
// (7, 5, 'neigh_op_bot_6')
// (8, 3, 'neigh_op_tnl_6')
// (8, 4, 'neigh_op_lft_6')
// (8, 5, 'neigh_op_bnl_6')

reg n306 = 0;
// (6, 3, 'neigh_op_tnr_7')
// (6, 4, 'neigh_op_rgt_7')
// (6, 5, 'neigh_op_bnr_7')
// (7, 3, 'local_g0_7')
// (7, 3, 'lutff_2/in_1')
// (7, 3, 'neigh_op_top_7')
// (7, 4, 'local_g2_7')
// (7, 4, 'lutff_0/in_1')
// (7, 4, 'lutff_7/out')
// (7, 5, 'neigh_op_bot_7')
// (8, 3, 'neigh_op_tnl_7')
// (8, 4, 'neigh_op_lft_7')
// (8, 5, 'neigh_op_bnl_7')

wire n307;
// (6, 4, 'neigh_op_tnr_0')
// (6, 5, 'neigh_op_rgt_0')
// (6, 6, 'neigh_op_bnr_0')
// (7, 1, 'sp12_v_t_23')
// (7, 2, 'sp12_v_b_23')
// (7, 3, 'sp12_v_b_20')
// (7, 3, 'sp4_r_v_b_41')
// (7, 4, 'neigh_op_top_0')
// (7, 4, 'sp12_v_b_19')
// (7, 4, 'sp4_r_v_b_28')
// (7, 5, 'lutff_0/out')
// (7, 5, 'sp12_v_b_16')
// (7, 5, 'sp4_r_v_b_17')
// (7, 6, 'neigh_op_bot_0')
// (7, 6, 'sp12_v_b_15')
// (7, 6, 'sp4_r_v_b_4')
// (7, 7, 'sp12_v_b_12')
// (7, 7, 'sp4_r_v_b_42')
// (7, 8, 'sp12_v_b_11')
// (7, 8, 'sp4_r_v_b_31')
// (7, 9, 'local_g2_0')
// (7, 9, 'local_g3_0')
// (7, 9, 'lutff_5/in_3')
// (7, 9, 'lutff_6/in_3')
// (7, 9, 'sp12_v_b_8')
// (7, 9, 'sp4_r_v_b_18')
// (7, 10, 'sp12_v_b_7')
// (7, 10, 'sp4_r_v_b_7')
// (7, 11, 'sp12_v_b_4')
// (7, 12, 'sp12_v_b_3')
// (7, 13, 'sp12_v_b_0')
// (8, 2, 'sp4_v_t_41')
// (8, 3, 'sp4_v_b_41')
// (8, 4, 'neigh_op_tnl_0')
// (8, 4, 'sp4_v_b_28')
// (8, 5, 'neigh_op_lft_0')
// (8, 5, 'sp4_v_b_17')
// (8, 6, 'neigh_op_bnl_0')
// (8, 6, 'sp4_v_b_4')
// (8, 6, 'sp4_v_t_42')
// (8, 7, 'sp4_v_b_42')
// (8, 8, 'sp4_v_b_31')
// (8, 9, 'local_g0_2')
// (8, 9, 'lutff_0/in_2')
// (8, 9, 'lutff_1/in_3')
// (8, 9, 'sp4_v_b_18')
// (8, 10, 'sp4_v_b_7')

reg n308 = 0;
// (6, 4, 'neigh_op_tnr_2')
// (6, 5, 'local_g3_2')
// (6, 5, 'lutff_1/in_0')
// (6, 5, 'neigh_op_rgt_2')
// (6, 6, 'neigh_op_bnr_2')
// (7, 4, 'neigh_op_top_2')
// (7, 5, 'lutff_2/out')
// (7, 6, 'neigh_op_bot_2')
// (8, 4, 'neigh_op_tnl_2')
// (8, 5, 'neigh_op_lft_2')
// (8, 6, 'neigh_op_bnl_2')

reg n309 = 0;
// (6, 4, 'neigh_op_tnr_4')
// (6, 5, 'neigh_op_rgt_4')
// (6, 6, 'neigh_op_bnr_4')
// (7, 4, 'neigh_op_top_4')
// (7, 5, 'local_g3_4')
// (7, 5, 'lutff_1/in_0')
// (7, 5, 'lutff_2/in_1')
// (7, 5, 'lutff_4/out')
// (7, 6, 'neigh_op_bot_4')
// (8, 4, 'neigh_op_tnl_4')
// (8, 5, 'neigh_op_lft_4')
// (8, 6, 'neigh_op_bnl_4')

reg n310 = 0;
// (6, 4, 'neigh_op_tnr_5')
// (6, 5, 'neigh_op_rgt_5')
// (6, 6, 'neigh_op_bnr_5')
// (7, 4, 'neigh_op_top_5')
// (7, 5, 'local_g1_5')
// (7, 5, 'lutff_4/in_0')
// (7, 5, 'lutff_5/out')
// (7, 6, 'neigh_op_bot_5')
// (8, 4, 'neigh_op_tnl_5')
// (8, 5, 'neigh_op_lft_5')
// (8, 6, 'neigh_op_bnl_5')

reg n311 = 0;
// (6, 4, 'neigh_op_tnr_6')
// (6, 5, 'neigh_op_rgt_6')
// (6, 6, 'neigh_op_bnr_6')
// (7, 4, 'neigh_op_top_6')
// (7, 5, 'local_g1_6')
// (7, 5, 'lutff_6/out')
// (7, 5, 'lutff_7/in_0')
// (7, 6, 'neigh_op_bot_6')
// (8, 4, 'neigh_op_tnl_6')
// (8, 5, 'neigh_op_lft_6')
// (8, 6, 'neigh_op_bnl_6')

reg n312 = 0;
// (6, 4, 'neigh_op_tnr_7')
// (6, 5, 'neigh_op_rgt_7')
// (6, 6, 'neigh_op_bnr_7')
// (7, 4, 'neigh_op_top_7')
// (7, 5, 'local_g0_7')
// (7, 5, 'lutff_5/in_0')
// (7, 5, 'lutff_7/out')
// (7, 6, 'neigh_op_bot_7')
// (8, 4, 'neigh_op_tnl_7')
// (8, 5, 'neigh_op_lft_7')
// (8, 6, 'neigh_op_bnl_7')

reg n313 = 0;
// (6, 4, 'sp12_h_r_1')
// (7, 4, 'sp12_h_r_2')
// (8, 3, 'neigh_op_tnr_7')
// (8, 4, 'neigh_op_rgt_7')
// (8, 4, 'sp12_h_r_5')
// (8, 5, 'neigh_op_bnr_7')
// (9, 3, 'neigh_op_top_7')
// (9, 4, 'local_g1_7')
// (9, 4, 'lutff_0/in_2')
// (9, 4, 'lutff_7/out')
// (9, 4, 'sp12_h_r_6')
// (9, 4, 'sp4_r_v_b_47')
// (9, 5, 'neigh_op_bot_7')
// (9, 5, 'sp4_r_v_b_34')
// (9, 6, 'sp4_r_v_b_23')
// (9, 7, 'sp4_r_v_b_10')
// (10, 3, 'neigh_op_tnl_7')
// (10, 3, 'sp4_h_r_3')
// (10, 3, 'sp4_v_t_47')
// (10, 4, 'neigh_op_lft_7')
// (10, 4, 'sp12_h_r_9')
// (10, 4, 'sp4_v_b_47')
// (10, 5, 'neigh_op_bnl_7')
// (10, 5, 'sp4_v_b_34')
// (10, 6, 'sp4_v_b_23')
// (10, 7, 'sp4_v_b_10')
// (11, 3, 'local_g0_6')
// (11, 3, 'lutff_1/in_3')
// (11, 3, 'sp4_h_r_14')
// (11, 4, 'local_g0_2')
// (11, 4, 'lutff_3/in_3')
// (11, 4, 'sp12_h_r_10')
// (12, 3, 'sp4_h_r_27')
// (12, 4, 'sp12_h_r_13')
// (13, 3, 'span4_horz_27')
// (13, 4, 'span12_horz_13')

reg n314 = 0;
// (6, 4, 'sp4_r_v_b_44')
// (6, 5, 'neigh_op_tnr_2')
// (6, 5, 'sp4_r_v_b_33')
// (6, 6, 'neigh_op_rgt_2')
// (6, 6, 'sp4_r_v_b_20')
// (6, 7, 'neigh_op_bnr_2')
// (6, 7, 'sp4_r_v_b_9')
// (7, 3, 'sp4_v_t_44')
// (7, 4, 'sp4_v_b_44')
// (7, 5, 'neigh_op_top_2')
// (7, 5, 'sp4_v_b_33')
// (7, 6, 'local_g0_2')
// (7, 6, 'lutff_2/out')
// (7, 6, 'lutff_4/in_0')
// (7, 6, 'sp4_v_b_20')
// (7, 7, 'local_g0_1')
// (7, 7, 'local_g0_2')
// (7, 7, 'lutff_1/in_1')
// (7, 7, 'lutff_4/in_2')
// (7, 7, 'lutff_7/in_0')
// (7, 7, 'neigh_op_bot_2')
// (7, 7, 'sp4_v_b_9')
// (8, 5, 'neigh_op_tnl_2')
// (8, 6, 'neigh_op_lft_2')
// (8, 7, 'neigh_op_bnl_2')

reg n315 = 0;
// (6, 5, 'neigh_op_tnr_0')
// (6, 6, 'neigh_op_rgt_0')
// (6, 7, 'neigh_op_bnr_0')
// (7, 5, 'neigh_op_top_0')
// (7, 6, 'local_g1_0')
// (7, 6, 'lutff_0/out')
// (7, 6, 'lutff_5/in_0')
// (7, 7, 'neigh_op_bot_0')
// (8, 5, 'neigh_op_tnl_0')
// (8, 6, 'neigh_op_lft_0')
// (8, 7, 'neigh_op_bnl_0')

reg n316 = 0;
// (6, 5, 'neigh_op_tnr_1')
// (6, 6, 'neigh_op_rgt_1')
// (6, 7, 'neigh_op_bnr_1')
// (7, 5, 'neigh_op_top_1')
// (7, 6, 'local_g0_1')
// (7, 6, 'lutff_1/out')
// (7, 6, 'lutff_7/in_0')
// (7, 7, 'neigh_op_bot_1')
// (8, 5, 'neigh_op_tnl_1')
// (8, 6, 'neigh_op_lft_1')
// (8, 7, 'neigh_op_bnl_1')

reg n317 = 0;
// (6, 5, 'neigh_op_tnr_3')
// (6, 6, 'neigh_op_rgt_3')
// (6, 7, 'neigh_op_bnr_3')
// (7, 5, 'neigh_op_top_3')
// (7, 6, 'local_g1_3')
// (7, 6, 'lutff_0/in_0')
// (7, 6, 'lutff_3/out')
// (7, 7, 'neigh_op_bot_3')
// (8, 5, 'neigh_op_tnl_3')
// (8, 6, 'neigh_op_lft_3')
// (8, 7, 'neigh_op_bnl_3')

reg n318 = 0;
// (6, 5, 'neigh_op_tnr_4')
// (6, 6, 'neigh_op_rgt_4')
// (6, 7, 'neigh_op_bnr_4')
// (7, 5, 'neigh_op_top_4')
// (7, 6, 'local_g1_4')
// (7, 6, 'lutff_1/in_0')
// (7, 6, 'lutff_4/out')
// (7, 7, 'neigh_op_bot_4')
// (8, 5, 'neigh_op_tnl_4')
// (8, 6, 'neigh_op_lft_4')
// (8, 7, 'neigh_op_bnl_4')

reg n319 = 0;
// (6, 5, 'neigh_op_tnr_6')
// (6, 6, 'neigh_op_rgt_6')
// (6, 7, 'neigh_op_bnr_6')
// (7, 5, 'neigh_op_top_6')
// (7, 6, 'local_g1_6')
// (7, 6, 'lutff_3/in_0')
// (7, 6, 'lutff_6/out')
// (7, 7, 'neigh_op_bot_6')
// (8, 5, 'neigh_op_tnl_6')
// (8, 6, 'neigh_op_lft_6')
// (8, 7, 'neigh_op_bnl_6')

reg n320 = 0;
// (6, 5, 'neigh_op_tnr_7')
// (6, 6, 'neigh_op_rgt_7')
// (6, 7, 'neigh_op_bnr_7')
// (7, 5, 'neigh_op_top_7')
// (7, 6, 'local_g1_7')
// (7, 6, 'lutff_2/in_0')
// (7, 6, 'lutff_7/out')
// (7, 7, 'neigh_op_bot_7')
// (8, 5, 'neigh_op_tnl_7')
// (8, 6, 'neigh_op_lft_7')
// (8, 7, 'neigh_op_bnl_7')

wire n321;
// (6, 5, 'sp4_r_v_b_47')
// (6, 6, 'sp4_r_v_b_34')
// (6, 7, 'sp4_r_v_b_23')
// (6, 8, 'sp4_r_v_b_10')
// (6, 11, 'neigh_op_tnr_6')
// (6, 12, 'neigh_op_rgt_6')
// (6, 13, 'neigh_op_bnr_6')
// (7, 4, 'sp4_v_t_47')
// (7, 5, 'sp4_v_b_47')
// (7, 6, 'sp12_v_t_23')
// (7, 6, 'sp4_v_b_34')
// (7, 7, 'sp12_v_b_23')
// (7, 7, 'sp4_v_b_23')
// (7, 8, 'sp12_v_b_20')
// (7, 8, 'sp4_h_r_4')
// (7, 8, 'sp4_v_b_10')
// (7, 9, 'local_g2_3')
// (7, 9, 'lutff_7/in_2')
// (7, 9, 'sp12_v_b_19')
// (7, 10, 'sp12_v_b_16')
// (7, 11, 'neigh_op_top_6')
// (7, 11, 'sp12_v_b_15')
// (7, 12, 'lutff_6/out')
// (7, 12, 'sp12_v_b_12')
// (7, 13, 'neigh_op_bot_6')
// (7, 13, 'sp12_v_b_11')
// (7, 14, 'sp12_v_b_8')
// (7, 15, 'sp12_v_b_7')
// (7, 16, 'sp12_v_b_4')
// (7, 17, 'span12_vert_3')
// (8, 8, 'local_g0_1')
// (8, 8, 'lutff_4/in_1')
// (8, 8, 'lutff_6/in_1')
// (8, 8, 'sp4_h_r_17')
// (8, 11, 'neigh_op_tnl_6')
// (8, 12, 'neigh_op_lft_6')
// (8, 13, 'neigh_op_bnl_6')
// (9, 8, 'sp4_h_r_28')
// (10, 8, 'sp4_h_r_41')
// (11, 8, 'sp4_h_l_41')

wire n322;
// (6, 6, 'neigh_op_tnr_0')
// (6, 6, 'sp4_r_v_b_45')
// (6, 7, 'neigh_op_rgt_0')
// (6, 7, 'sp4_r_v_b_32')
// (6, 8, 'neigh_op_bnr_0')
// (6, 8, 'sp4_r_v_b_21')
// (6, 9, 'sp4_r_v_b_8')
// (7, 5, 'sp4_v_t_45')
// (7, 6, 'neigh_op_top_0')
// (7, 6, 'sp4_v_b_45')
// (7, 7, 'lutff_0/out')
// (7, 7, 'sp4_v_b_32')
// (7, 8, 'neigh_op_bot_0')
// (7, 8, 'sp4_v_b_21')
// (7, 9, 'local_g1_0')
// (7, 9, 'lutff_5/in_0')
// (7, 9, 'sp4_v_b_8')
// (8, 6, 'neigh_op_tnl_0')
// (8, 7, 'neigh_op_lft_0')
// (8, 8, 'neigh_op_bnl_0')

wire n323;
// (6, 6, 'neigh_op_tnr_1')
// (6, 7, 'neigh_op_rgt_1')
// (6, 8, 'neigh_op_bnr_1')
// (7, 6, 'neigh_op_top_1')
// (7, 7, 'local_g2_1')
// (7, 7, 'lutff_0/in_3')
// (7, 7, 'lutff_1/out')
// (7, 8, 'neigh_op_bot_1')
// (8, 6, 'neigh_op_tnl_1')
// (8, 7, 'neigh_op_lft_1')
// (8, 8, 'neigh_op_bnl_1')

reg n324 = 0;
// (6, 6, 'neigh_op_tnr_2')
// (6, 7, 'neigh_op_rgt_2')
// (6, 8, 'neigh_op_bnr_2')
// (7, 6, 'neigh_op_top_2')
// (7, 7, 'local_g1_2')
// (7, 7, 'lutff_2/out')
// (7, 7, 'lutff_3/in_0')
// (7, 8, 'neigh_op_bot_2')
// (8, 6, 'neigh_op_tnl_2')
// (8, 7, 'neigh_op_lft_2')
// (8, 8, 'neigh_op_bnl_2')

reg n325 = 0;
// (6, 6, 'neigh_op_tnr_3')
// (6, 7, 'neigh_op_rgt_3')
// (6, 8, 'neigh_op_bnr_3')
// (7, 6, 'neigh_op_top_3')
// (7, 7, 'local_g1_3')
// (7, 7, 'lutff_3/out')
// (7, 7, 'lutff_6/in_0')
// (7, 8, 'neigh_op_bot_3')
// (8, 6, 'neigh_op_tnl_3')
// (8, 7, 'neigh_op_lft_3')
// (8, 8, 'neigh_op_bnl_3')

reg n326 = 0;
// (6, 6, 'neigh_op_tnr_4')
// (6, 7, 'neigh_op_rgt_4')
// (6, 8, 'neigh_op_bnr_4')
// (7, 6, 'neigh_op_top_4')
// (7, 7, 'local_g2_4')
// (7, 7, 'lutff_2/in_0')
// (7, 7, 'lutff_4/out')
// (7, 8, 'neigh_op_bot_4')
// (8, 6, 'neigh_op_tnl_4')
// (8, 7, 'neigh_op_lft_4')
// (8, 8, 'neigh_op_bnl_4')

reg n327 = 0;
// (6, 6, 'neigh_op_tnr_5')
// (6, 7, 'neigh_op_rgt_5')
// (6, 8, 'neigh_op_bnr_5')
// (7, 6, 'neigh_op_top_5')
// (7, 7, 'lutff_5/out')
// (7, 8, 'local_g0_5')
// (7, 8, 'lutff_1/in_0')
// (7, 8, 'neigh_op_bot_5')
// (8, 6, 'neigh_op_tnl_5')
// (8, 7, 'neigh_op_lft_5')
// (8, 8, 'neigh_op_bnl_5')

reg n328 = 0;
// (6, 6, 'neigh_op_tnr_6')
// (6, 7, 'neigh_op_rgt_6')
// (6, 8, 'neigh_op_bnr_6')
// (7, 6, 'neigh_op_top_6')
// (7, 7, 'local_g0_6')
// (7, 7, 'local_g1_6')
// (7, 7, 'lutff_1/in_0')
// (7, 7, 'lutff_6/out')
// (7, 7, 'lutff_7/in_1')
// (7, 8, 'neigh_op_bot_6')
// (8, 6, 'neigh_op_tnl_6')
// (8, 7, 'neigh_op_lft_6')
// (8, 8, 'neigh_op_bnl_6')

reg n329 = 0;
// (6, 6, 'neigh_op_tnr_7')
// (6, 7, 'neigh_op_rgt_7')
// (6, 8, 'neigh_op_bnr_7')
// (7, 6, 'neigh_op_top_7')
// (7, 7, 'local_g0_7')
// (7, 7, 'lutff_5/in_0')
// (7, 7, 'lutff_7/out')
// (7, 8, 'neigh_op_bot_7')
// (8, 6, 'neigh_op_tnl_7')
// (8, 7, 'neigh_op_lft_7')
// (8, 8, 'neigh_op_bnl_7')

reg n330 = 0;
// (6, 7, 'neigh_op_tnr_1')
// (6, 8, 'neigh_op_rgt_1')
// (6, 9, 'neigh_op_bnr_1')
// (7, 7, 'neigh_op_top_1')
// (7, 8, 'local_g0_1')
// (7, 8, 'lutff_1/out')
// (7, 8, 'lutff_5/in_0')
// (7, 9, 'neigh_op_bot_1')
// (8, 7, 'neigh_op_tnl_1')
// (8, 8, 'neigh_op_lft_1')
// (8, 9, 'neigh_op_bnl_1')

reg n331 = 0;
// (6, 7, 'neigh_op_tnr_5')
// (6, 8, 'neigh_op_rgt_5')
// (6, 9, 'neigh_op_bnr_5')
// (7, 5, 'sp4_r_v_b_46')
// (7, 6, 'local_g2_3')
// (7, 6, 'lutff_4/in_1')
// (7, 6, 'sp4_r_v_b_35')
// (7, 7, 'local_g1_5')
// (7, 7, 'lutff_0/in_0')
// (7, 7, 'neigh_op_top_5')
// (7, 7, 'sp4_r_v_b_22')
// (7, 8, 'lutff_5/out')
// (7, 8, 'sp4_r_v_b_11')
// (7, 9, 'neigh_op_bot_5')
// (8, 4, 'sp4_v_t_46')
// (8, 5, 'sp4_v_b_46')
// (8, 6, 'sp4_v_b_35')
// (8, 7, 'neigh_op_tnl_5')
// (8, 7, 'sp4_v_b_22')
// (8, 8, 'neigh_op_lft_5')
// (8, 8, 'sp4_v_b_11')
// (8, 9, 'neigh_op_bnl_5')

reg n332 = 0;
// (6, 7, 'sp4_h_r_5')
// (7, 7, 'sp4_h_r_16')
// (8, 6, 'neigh_op_tnr_4')
// (8, 7, 'neigh_op_rgt_4')
// (8, 7, 'sp4_h_r_29')
// (8, 8, 'neigh_op_bnr_4')
// (9, 6, 'neigh_op_top_4')
// (9, 7, 'local_g2_0')
// (9, 7, 'local_g3_0')
// (9, 7, 'lutff_2/in_1')
// (9, 7, 'lutff_3/in_1')
// (9, 7, 'lutff_4/out')
// (9, 7, 'sp4_h_r_40')
// (9, 8, 'neigh_op_bot_4')
// (10, 6, 'neigh_op_tnl_4')
// (10, 7, 'neigh_op_lft_4')
// (10, 7, 'sp4_h_l_40')
// (10, 8, 'neigh_op_bnl_4')

wire n333;
// (6, 8, 'local_g2_4')
// (6, 8, 'lutff_7/in_3')
// (6, 8, 'neigh_op_tnr_4')
// (6, 9, 'neigh_op_rgt_4')
// (6, 10, 'neigh_op_bnr_4')
// (7, 8, 'neigh_op_top_4')
// (7, 9, 'lutff_4/out')
// (7, 10, 'neigh_op_bot_4')
// (8, 8, 'neigh_op_tnl_4')
// (8, 9, 'neigh_op_lft_4')
// (8, 10, 'neigh_op_bnl_4')

wire n334;
// (6, 8, 'neigh_op_tnr_6')
// (6, 9, 'neigh_op_rgt_6')
// (6, 9, 'sp4_h_r_1')
// (6, 10, 'neigh_op_bnr_6')
// (7, 7, 'sp4_r_v_b_37')
// (7, 8, 'neigh_op_top_6')
// (7, 8, 'sp4_r_v_b_24')
// (7, 9, 'lutff_6/out')
// (7, 9, 'sp4_h_r_12')
// (7, 9, 'sp4_r_v_b_13')
// (7, 10, 'neigh_op_bot_6')
// (7, 10, 'sp4_r_v_b_0')
// (8, 6, 'sp4_v_t_37')
// (8, 7, 'sp4_v_b_37')
// (8, 8, 'neigh_op_tnl_6')
// (8, 8, 'sp4_v_b_24')
// (8, 9, 'neigh_op_lft_6')
// (8, 9, 'sp4_h_r_25')
// (8, 9, 'sp4_v_b_13')
// (8, 10, 'local_g2_6')
// (8, 10, 'local_g3_6')
// (8, 10, 'lutff_0/in_3')
// (8, 10, 'lutff_1/in_1')
// (8, 10, 'lutff_2/in_2')
// (8, 10, 'lutff_3/in_2')
// (8, 10, 'neigh_op_bnl_6')
// (8, 10, 'sp4_h_r_6')
// (8, 10, 'sp4_v_b_0')
// (9, 9, 'sp4_h_r_36')
// (9, 10, 'local_g0_3')
// (9, 10, 'local_g2_4')
// (9, 10, 'lutff_0/in_0')
// (9, 10, 'lutff_1/in_0')
// (9, 10, 'lutff_3/in_1')
// (9, 10, 'lutff_4/in_0')
// (9, 10, 'lutff_5/in_2')
// (9, 10, 'sp4_h_r_19')
// (9, 10, 'sp4_r_v_b_36')
// (9, 11, 'sp4_r_v_b_25')
// (9, 12, 'sp4_r_v_b_12')
// (9, 13, 'sp4_r_v_b_1')
// (10, 9, 'sp4_h_l_36')
// (10, 9, 'sp4_v_t_36')
// (10, 10, 'sp4_h_r_30')
// (10, 10, 'sp4_v_b_36')
// (10, 11, 'sp4_v_b_25')
// (10, 12, 'sp4_v_b_12')
// (10, 13, 'sp4_v_b_1')
// (11, 10, 'sp4_h_r_43')
// (12, 10, 'sp4_h_l_43')

reg n335 = 0;
// (6, 8, 'neigh_op_tnr_7')
// (6, 9, 'local_g3_7')
// (6, 9, 'lutff_6/in_0')
// (6, 9, 'neigh_op_rgt_7')
// (6, 10, 'neigh_op_bnr_7')
// (7, 8, 'neigh_op_top_7')
// (7, 9, 'lutff_7/out')
// (7, 10, 'neigh_op_bot_7')
// (8, 8, 'neigh_op_tnl_7')
// (8, 9, 'neigh_op_lft_7')
// (8, 10, 'neigh_op_bnl_7')

wire n336;
// (6, 8, 'sp4_r_v_b_46')
// (6, 9, 'sp4_r_v_b_35')
// (6, 10, 'sp4_r_v_b_22')
// (6, 11, 'sp4_r_v_b_11')
// (7, 7, 'sp4_v_t_46')
// (7, 8, 'sp4_v_b_46')
// (7, 9, 'sp4_v_b_35')
// (7, 10, 'sp4_v_b_22')
// (7, 11, 'local_g0_3')
// (7, 11, 'local_g1_3')
// (7, 11, 'lutff_0/in_2')
// (7, 11, 'lutff_1/in_0')
// (7, 11, 'lutff_2/in_2')
// (7, 11, 'lutff_3/in_3')
// (7, 11, 'lutff_4/in_3')
// (7, 11, 'lutff_6/in_1')
// (7, 11, 'sp4_h_r_6')
// (7, 11, 'sp4_v_b_11')
// (8, 10, 'neigh_op_tnr_7')
// (8, 11, 'local_g2_7')
// (8, 11, 'local_g3_7')
// (8, 11, 'lutff_6/in_1')
// (8, 11, 'lutff_7/in_1')
// (8, 11, 'neigh_op_rgt_7')
// (8, 11, 'sp4_h_r_19')
// (8, 12, 'neigh_op_bnr_7')
// (9, 10, 'neigh_op_top_7')
// (9, 11, 'lutff_7/out')
// (9, 11, 'sp4_h_r_30')
// (9, 12, 'neigh_op_bot_7')
// (10, 10, 'neigh_op_tnl_7')
// (10, 11, 'neigh_op_lft_7')
// (10, 11, 'sp4_h_r_43')
// (10, 12, 'neigh_op_bnl_7')
// (11, 11, 'sp4_h_l_43')

wire n337;
// (6, 9, 'neigh_op_tnr_1')
// (6, 10, 'neigh_op_rgt_1')
// (6, 11, 'neigh_op_bnr_1')
// (7, 9, 'local_g0_1')
// (7, 9, 'local_g1_1')
// (7, 9, 'lutff_0/in_2')
// (7, 9, 'lutff_3/in_2')
// (7, 9, 'neigh_op_top_1')
// (7, 10, 'lutff_1/out')
// (7, 11, 'neigh_op_bot_1')
// (8, 9, 'local_g3_1')
// (8, 9, 'lutff_7/in_1')
// (8, 9, 'neigh_op_tnl_1')
// (8, 10, 'neigh_op_lft_1')
// (8, 11, 'neigh_op_bnl_1')

wire n338;
// (6, 9, 'neigh_op_tnr_2')
// (6, 10, 'neigh_op_rgt_2')
// (6, 11, 'neigh_op_bnr_2')
// (7, 9, 'local_g1_2')
// (7, 9, 'lutff_1/in_2')
// (7, 9, 'neigh_op_top_2')
// (7, 10, 'lutff_2/out')
// (7, 11, 'neigh_op_bot_2')
// (8, 9, 'local_g2_2')
// (8, 9, 'local_g3_2')
// (8, 9, 'lutff_3/in_2')
// (8, 9, 'lutff_5/in_0')
// (8, 9, 'lutff_6/in_0')
// (8, 9, 'neigh_op_tnl_2')
// (8, 10, 'neigh_op_lft_2')
// (8, 11, 'neigh_op_bnl_2')

wire n339;
// (6, 9, 'neigh_op_tnr_3')
// (6, 10, 'neigh_op_rgt_3')
// (6, 11, 'neigh_op_bnr_3')
// (7, 9, 'neigh_op_top_3')
// (7, 10, 'local_g0_3')
// (7, 10, 'lutff_3/out')
// (7, 10, 'lutff_6/in_3')
// (7, 11, 'neigh_op_bot_3')
// (8, 9, 'neigh_op_tnl_3')
// (8, 10, 'neigh_op_lft_3')
// (8, 11, 'neigh_op_bnl_3')

wire n340;
// (6, 9, 'neigh_op_tnr_4')
// (6, 10, 'neigh_op_rgt_4')
// (6, 11, 'neigh_op_bnr_4')
// (7, 9, 'local_g1_4')
// (7, 9, 'lutff_4/in_3')
// (7, 9, 'neigh_op_top_4')
// (7, 10, 'local_g3_1')
// (7, 10, 'lutff_4/out')
// (7, 10, 'lutff_6/in_2')
// (7, 10, 'lutff_7/in_3')
// (7, 10, 'sp4_r_v_b_41')
// (7, 11, 'neigh_op_bot_4')
// (7, 11, 'sp4_r_v_b_28')
// (7, 12, 'sp4_r_v_b_17')
// (7, 13, 'sp4_r_v_b_4')
// (8, 9, 'neigh_op_tnl_4')
// (8, 9, 'sp4_v_t_41')
// (8, 10, 'neigh_op_lft_4')
// (8, 10, 'sp4_v_b_41')
// (8, 11, 'neigh_op_bnl_4')
// (8, 11, 'sp4_v_b_28')
// (8, 12, 'sp4_v_b_17')
// (8, 13, 'sp4_v_b_4')

wire n341;
// (6, 9, 'neigh_op_tnr_5')
// (6, 10, 'neigh_op_rgt_5')
// (6, 11, 'neigh_op_bnr_5')
// (7, 9, 'neigh_op_top_5')
// (7, 10, 'lutff_5/out')
// (7, 11, 'neigh_op_bot_5')
// (8, 9, 'local_g3_5')
// (8, 9, 'lutff_5/in_3')
// (8, 9, 'neigh_op_tnl_5')
// (8, 10, 'neigh_op_lft_5')
// (8, 11, 'neigh_op_bnl_5')

wire n342;
// (6, 10, 'neigh_op_tnr_0')
// (6, 11, 'neigh_op_rgt_0')
// (6, 12, 'neigh_op_bnr_0')
// (7, 10, 'local_g0_0')
// (7, 10, 'local_g1_0')
// (7, 10, 'lutff_3/in_0')
// (7, 10, 'lutff_4/in_0')
// (7, 10, 'neigh_op_top_0')
// (7, 11, 'lutff_0/out')
// (7, 12, 'neigh_op_bot_0')
// (8, 10, 'neigh_op_tnl_0')
// (8, 11, 'neigh_op_lft_0')
// (8, 12, 'neigh_op_bnl_0')

wire n343;
// (6, 10, 'neigh_op_tnr_1')
// (6, 11, 'neigh_op_rgt_1')
// (6, 12, 'neigh_op_bnr_1')
// (7, 10, 'local_g1_1')
// (7, 10, 'lutff_2/in_0')
// (7, 10, 'lutff_5/in_1')
// (7, 10, 'neigh_op_top_1')
// (7, 11, 'lutff_1/out')
// (7, 12, 'neigh_op_bot_1')
// (8, 10, 'neigh_op_tnl_1')
// (8, 11, 'neigh_op_lft_1')
// (8, 12, 'neigh_op_bnl_1')

wire n344;
// (6, 10, 'neigh_op_tnr_2')
// (6, 11, 'neigh_op_rgt_2')
// (6, 12, 'neigh_op_bnr_2')
// (7, 10, 'neigh_op_top_2')
// (7, 11, 'lutff_2/out')
// (7, 12, 'neigh_op_bot_2')
// (8, 10, 'neigh_op_tnl_2')
// (8, 11, 'local_g0_2')
// (8, 11, 'local_g1_2')
// (8, 11, 'lutff_0/in_0')
// (8, 11, 'lutff_1/in_0')
// (8, 11, 'lutff_2/in_0')
// (8, 11, 'lutff_4/in_0')
// (8, 11, 'neigh_op_lft_2')
// (8, 12, 'neigh_op_bnl_2')

wire n345;
// (6, 10, 'neigh_op_tnr_3')
// (6, 11, 'neigh_op_rgt_3')
// (6, 12, 'neigh_op_bnr_3')
// (7, 10, 'neigh_op_top_3')
// (7, 11, 'lutff_3/out')
// (7, 12, 'neigh_op_bot_3')
// (8, 10, 'local_g2_3')
// (8, 10, 'local_g3_3')
// (8, 10, 'lutff_4/in_0')
// (8, 10, 'lutff_5/in_0')
// (8, 10, 'neigh_op_tnl_3')
// (8, 11, 'neigh_op_lft_3')
// (8, 12, 'neigh_op_bnl_3')

wire n346;
// (6, 10, 'neigh_op_tnr_4')
// (6, 11, 'neigh_op_rgt_4')
// (6, 12, 'neigh_op_bnr_4')
// (7, 10, 'local_g0_4')
// (7, 10, 'local_g1_4')
// (7, 10, 'lutff_2/in_2')
// (7, 10, 'lutff_3/in_2')
// (7, 10, 'lutff_4/in_2')
// (7, 10, 'lutff_5/in_2')
// (7, 10, 'neigh_op_top_4')
// (7, 11, 'lutff_4/out')
// (7, 12, 'neigh_op_bot_4')
// (8, 10, 'neigh_op_tnl_4')
// (8, 11, 'neigh_op_lft_4')
// (8, 12, 'neigh_op_bnl_4')

wire n347;
// (6, 10, 'neigh_op_tnr_6')
// (6, 11, 'neigh_op_rgt_6')
// (6, 12, 'neigh_op_bnr_6')
// (7, 10, 'neigh_op_top_6')
// (7, 11, 'lutff_6/out')
// (7, 12, 'neigh_op_bot_6')
// (8, 10, 'neigh_op_tnl_6')
// (8, 11, 'local_g0_6')
// (8, 11, 'local_g1_6')
// (8, 11, 'lutff_0/in_1')
// (8, 11, 'lutff_1/in_1')
// (8, 11, 'lutff_2/in_1')
// (8, 11, 'lutff_4/in_1')
// (8, 11, 'neigh_op_lft_6')
// (8, 12, 'neigh_op_bnl_6')

wire n348;
// (6, 10, 'sp4_h_r_3')
// (7, 10, 'local_g0_6')
// (7, 10, 'local_g1_6')
// (7, 10, 'lutff_2/in_1')
// (7, 10, 'lutff_3/in_3')
// (7, 10, 'sp4_h_r_14')
// (8, 8, 'sp4_r_v_b_46')
// (8, 9, 'neigh_op_tnr_3')
// (8, 9, 'sp4_r_v_b_35')
// (8, 10, 'neigh_op_rgt_3')
// (8, 10, 'sp4_h_r_27')
// (8, 10, 'sp4_r_v_b_22')
// (8, 10, 'sp4_r_v_b_38')
// (8, 11, 'local_g2_3')
// (8, 11, 'lutff_5/in_2')
// (8, 11, 'neigh_op_bnr_3')
// (8, 11, 'sp4_r_v_b_11')
// (8, 11, 'sp4_r_v_b_27')
// (8, 12, 'sp4_r_v_b_14')
// (8, 13, 'sp4_r_v_b_3')
// (9, 7, 'sp4_v_t_46')
// (9, 8, 'sp4_v_b_46')
// (9, 9, 'neigh_op_top_3')
// (9, 9, 'sp4_v_b_35')
// (9, 9, 'sp4_v_t_38')
// (9, 10, 'lutff_3/out')
// (9, 10, 'sp4_h_r_38')
// (9, 10, 'sp4_v_b_22')
// (9, 10, 'sp4_v_b_38')
// (9, 11, 'local_g2_3')
// (9, 11, 'local_g3_3')
// (9, 11, 'lutff_0/in_1')
// (9, 11, 'lutff_3/in_1')
// (9, 11, 'neigh_op_bot_3')
// (9, 11, 'sp4_v_b_11')
// (9, 11, 'sp4_v_b_27')
// (9, 12, 'sp4_v_b_14')
// (9, 13, 'sp4_v_b_3')
// (10, 9, 'neigh_op_tnl_3')
// (10, 10, 'neigh_op_lft_3')
// (10, 10, 'sp4_h_l_38')
// (10, 11, 'neigh_op_bnl_3')

wire n349;
// (6, 11, 'neigh_op_tnr_0')
// (6, 12, 'neigh_op_rgt_0')
// (6, 13, 'neigh_op_bnr_0')
// (7, 11, 'neigh_op_top_0')
// (7, 12, 'local_g0_0')
// (7, 12, 'lutff_0/out')
// (7, 12, 'lutff_2/in_2')
// (7, 13, 'neigh_op_bot_0')
// (8, 11, 'neigh_op_tnl_0')
// (8, 12, 'neigh_op_lft_0')
// (8, 13, 'neigh_op_bnl_0')

wire n350;
// (6, 11, 'neigh_op_tnr_4')
// (6, 12, 'neigh_op_rgt_4')
// (6, 13, 'neigh_op_bnr_4')
// (7, 11, 'neigh_op_top_4')
// (7, 12, 'local_g2_4')
// (7, 12, 'lutff_4/out')
// (7, 12, 'lutff_6/in_2')
// (7, 13, 'neigh_op_bot_4')
// (8, 11, 'neigh_op_tnl_4')
// (8, 12, 'neigh_op_lft_4')
// (8, 13, 'neigh_op_bnl_4')

wire n351;
// (6, 11, 'neigh_op_tnr_7')
// (6, 12, 'neigh_op_rgt_7')
// (6, 13, 'neigh_op_bnr_7')
// (7, 11, 'neigh_op_top_7')
// (7, 12, 'local_g3_7')
// (7, 12, 'lutff_1/in_3')
// (7, 12, 'lutff_7/out')
// (7, 13, 'neigh_op_bot_7')
// (8, 11, 'neigh_op_tnl_7')
// (8, 12, 'neigh_op_lft_7')
// (8, 13, 'neigh_op_bnl_7')

wire n352;
// (6, 11, 'sp4_h_r_5')
// (7, 11, 'local_g0_0')
// (7, 11, 'local_g1_0')
// (7, 11, 'lutff_0/in_3')
// (7, 11, 'lutff_1/in_1')
// (7, 11, 'lutff_2/in_3')
// (7, 11, 'lutff_3/in_1')
// (7, 11, 'lutff_4/in_1')
// (7, 11, 'lutff_6/in_2')
// (7, 11, 'sp4_h_r_16')
// (8, 10, 'neigh_op_tnr_4')
// (8, 11, 'local_g2_4')
// (8, 11, 'lutff_6/in_0')
// (8, 11, 'lutff_7/in_3')
// (8, 11, 'neigh_op_rgt_4')
// (8, 11, 'sp4_h_r_29')
// (8, 12, 'neigh_op_bnr_4')
// (9, 10, 'neigh_op_top_4')
// (9, 11, 'lutff_4/out')
// (9, 11, 'sp4_h_r_40')
// (9, 12, 'neigh_op_bot_4')
// (10, 10, 'neigh_op_tnl_4')
// (10, 11, 'neigh_op_lft_4')
// (10, 11, 'sp4_h_l_40')
// (10, 12, 'neigh_op_bnl_4')

wire n353;
// (6, 11, 'sp4_h_r_7')
// (7, 11, 'local_g0_2')
// (7, 11, 'local_g1_2')
// (7, 11, 'lutff_0/in_1')
// (7, 11, 'lutff_1/in_2')
// (7, 11, 'lutff_2/in_1')
// (7, 11, 'lutff_3/in_0')
// (7, 11, 'lutff_4/in_2')
// (7, 11, 'lutff_6/in_3')
// (7, 11, 'sp4_h_r_18')
// (8, 10, 'neigh_op_tnr_5')
// (8, 11, 'local_g2_5')
// (8, 11, 'local_g3_5')
// (8, 11, 'lutff_6/in_2')
// (8, 11, 'lutff_7/in_0')
// (8, 11, 'neigh_op_rgt_5')
// (8, 11, 'sp4_h_r_31')
// (8, 12, 'neigh_op_bnr_5')
// (9, 10, 'neigh_op_top_5')
// (9, 11, 'lutff_5/out')
// (9, 11, 'sp4_h_r_42')
// (9, 12, 'neigh_op_bot_5')
// (10, 10, 'neigh_op_tnl_5')
// (10, 11, 'neigh_op_lft_5')
// (10, 11, 'sp4_h_l_42')
// (10, 12, 'neigh_op_bnl_5')

wire n354;
// (6, 11, 'sp4_r_v_b_43')
// (6, 12, 'local_g0_6')
// (6, 12, 'lutff_3/in_1')
// (6, 12, 'sp4_r_v_b_30')
// (6, 13, 'neigh_op_tnr_3')
// (6, 13, 'sp4_r_v_b_19')
// (6, 14, 'neigh_op_rgt_3')
// (6, 14, 'sp4_r_v_b_6')
// (6, 15, 'neigh_op_bnr_3')
// (7, 5, 'sp12_v_t_22')
// (7, 6, 'sp12_v_b_22')
// (7, 7, 'sp12_v_b_21')
// (7, 8, 'sp12_v_b_18')
// (7, 9, 'sp12_v_b_17')
// (7, 10, 'sp12_v_b_14')
// (7, 10, 'sp4_v_t_43')
// (7, 11, 'sp12_v_b_13')
// (7, 11, 'sp4_v_b_43')
// (7, 12, 'local_g2_2')
// (7, 12, 'local_g3_6')
// (7, 12, 'lutff_2/in_1')
// (7, 12, 'lutff_3/in_1')
// (7, 12, 'sp12_v_b_10')
// (7, 12, 'sp4_v_b_30')
// (7, 13, 'neigh_op_top_3')
// (7, 13, 'sp12_v_b_9')
// (7, 13, 'sp4_v_b_19')
// (7, 14, 'lutff_3/out')
// (7, 14, 'sp12_v_b_6')
// (7, 14, 'sp4_v_b_6')
// (7, 15, 'neigh_op_bot_3')
// (7, 15, 'sp12_v_b_5')
// (7, 16, 'sp12_v_b_2')
// (7, 17, 'span12_vert_1')
// (8, 13, 'neigh_op_tnl_3')
// (8, 14, 'neigh_op_lft_3')
// (8, 15, 'neigh_op_bnl_3')

wire n355;
// (6, 12, 'neigh_op_tnr_0')
// (6, 13, 'neigh_op_rgt_0')
// (6, 14, 'neigh_op_bnr_0')
// (7, 12, 'neigh_op_top_0')
// (7, 12, 'sp4_r_v_b_44')
// (7, 13, 'lutff_0/out')
// (7, 13, 'sp4_r_v_b_33')
// (7, 14, 'neigh_op_bot_0')
// (7, 14, 'sp4_r_v_b_20')
// (7, 15, 'sp4_r_v_b_9')
// (8, 11, 'sp4_v_t_44')
// (8, 12, 'neigh_op_tnl_0')
// (8, 12, 'sp4_v_b_44')
// (8, 13, 'local_g3_1')
// (8, 13, 'lutff_0/in_2')
// (8, 13, 'lutff_1/in_3')
// (8, 13, 'neigh_op_lft_0')
// (8, 13, 'sp4_v_b_33')
// (8, 14, 'neigh_op_bnl_0')
// (8, 14, 'sp4_v_b_20')
// (8, 15, 'sp4_v_b_9')

wire n356;
// (6, 12, 'neigh_op_tnr_1')
// (6, 13, 'neigh_op_rgt_1')
// (6, 14, 'neigh_op_bnr_1')
// (7, 12, 'neigh_op_top_1')
// (7, 13, 'lutff_1/out')
// (7, 14, 'neigh_op_bot_1')
// (8, 12, 'local_g3_1')
// (8, 12, 'lutff_3/in_3')
// (8, 12, 'lutff_7/in_3')
// (8, 12, 'neigh_op_tnl_1')
// (8, 13, 'local_g1_1')
// (8, 13, 'lutff_7/in_3')
// (8, 13, 'neigh_op_lft_1')
// (8, 14, 'neigh_op_bnl_1')

wire n357;
// (6, 12, 'neigh_op_tnr_2')
// (6, 13, 'neigh_op_rgt_2')
// (6, 13, 'sp4_r_v_b_36')
// (6, 14, 'local_g0_1')
// (6, 14, 'lutff_5/in_0')
// (6, 14, 'lutff_7/in_0')
// (6, 14, 'neigh_op_bnr_2')
// (6, 14, 'sp4_r_v_b_25')
// (6, 15, 'sp4_r_v_b_12')
// (6, 16, 'sp4_r_v_b_1')
// (7, 12, 'neigh_op_top_2')
// (7, 12, 'sp4_v_t_36')
// (7, 13, 'lutff_2/out')
// (7, 13, 'sp4_v_b_36')
// (7, 14, 'neigh_op_bot_2')
// (7, 14, 'sp4_v_b_25')
// (7, 15, 'sp4_v_b_12')
// (7, 16, 'sp4_v_b_1')
// (8, 12, 'neigh_op_tnl_2')
// (8, 13, 'neigh_op_lft_2')
// (8, 14, 'local_g2_2')
// (8, 14, 'local_g3_2')
// (8, 14, 'lutff_3/in_0')
// (8, 14, 'lutff_5/in_3')
// (8, 14, 'lutff_6/in_3')
// (8, 14, 'neigh_op_bnl_2')

wire n358;
// (6, 12, 'neigh_op_tnr_3')
// (6, 13, 'neigh_op_rgt_3')
// (6, 14, 'neigh_op_bnr_3')
// (7, 12, 'neigh_op_top_3')
// (7, 13, 'local_g0_3')
// (7, 13, 'lutff_3/out')
// (7, 13, 'lutff_6/in_3')
// (7, 14, 'neigh_op_bot_3')
// (8, 12, 'neigh_op_tnl_3')
// (8, 13, 'local_g1_3')
// (8, 13, 'lutff_6/in_2')
// (8, 13, 'neigh_op_lft_3')
// (8, 14, 'neigh_op_bnl_3')

wire n359;
// (6, 12, 'neigh_op_tnr_4')
// (6, 13, 'neigh_op_rgt_4')
// (6, 14, 'neigh_op_bnr_4')
// (7, 12, 'neigh_op_top_4')
// (7, 13, 'local_g0_4')
// (7, 13, 'local_g1_4')
// (7, 13, 'lutff_4/out')
// (7, 13, 'lutff_5/in_3')
// (7, 13, 'lutff_7/in_2')
// (7, 14, 'neigh_op_bot_4')
// (8, 12, 'neigh_op_tnl_4')
// (8, 13, 'neigh_op_lft_4')
// (8, 14, 'neigh_op_bnl_4')

wire n360;
// (6, 12, 'neigh_op_tnr_5')
// (6, 13, 'neigh_op_rgt_5')
// (6, 14, 'neigh_op_bnr_5')
// (7, 12, 'neigh_op_top_5')
// (7, 13, 'lutff_5/out')
// (7, 13, 'sp4_h_r_10')
// (7, 14, 'neigh_op_bot_5')
// (8, 12, 'neigh_op_tnl_5')
// (8, 13, 'local_g1_7')
// (8, 13, 'lutff_2/in_0')
// (8, 13, 'neigh_op_lft_5')
// (8, 13, 'sp4_h_r_23')
// (8, 14, 'neigh_op_bnl_5')
// (9, 13, 'sp4_h_r_34')
// (10, 13, 'sp4_h_r_47')
// (11, 13, 'sp4_h_l_47')

wire n361;
// (6, 12, 'neigh_op_tnr_6')
// (6, 13, 'neigh_op_rgt_6')
// (6, 14, 'neigh_op_bnr_6')
// (7, 12, 'local_g0_6')
// (7, 12, 'lutff_6/in_0')
// (7, 12, 'neigh_op_top_6')
// (7, 13, 'lutff_6/out')
// (7, 14, 'neigh_op_bot_6')
// (8, 12, 'neigh_op_tnl_6')
// (8, 13, 'neigh_op_lft_6')
// (8, 14, 'neigh_op_bnl_6')

wire n362;
// (6, 12, 'sp4_r_v_b_37')
// (6, 13, 'sp4_r_v_b_24')
// (6, 14, 'neigh_op_tnr_0')
// (6, 14, 'sp4_r_v_b_13')
// (6, 15, 'neigh_op_rgt_0')
// (6, 15, 'sp4_r_v_b_0')
// (6, 16, 'neigh_op_bnr_0')
// (7, 11, 'sp4_v_t_37')
// (7, 12, 'sp4_v_b_37')
// (7, 13, 'sp4_v_b_24')
// (7, 14, 'local_g1_0')
// (7, 14, 'local_g1_5')
// (7, 14, 'lutff_1/in_3')
// (7, 14, 'lutff_2/in_1')
// (7, 14, 'lutff_6/in_3')
// (7, 14, 'lutff_7/in_0')
// (7, 14, 'neigh_op_top_0')
// (7, 14, 'sp4_v_b_13')
// (7, 15, 'lutff_0/out')
// (7, 15, 'sp4_v_b_0')
// (7, 16, 'neigh_op_bot_0')
// (8, 14, 'local_g2_0')
// (8, 14, 'local_g3_0')
// (8, 14, 'lutff_0/in_1')
// (8, 14, 'lutff_1/in_3')
// (8, 14, 'lutff_2/in_3')
// (8, 14, 'neigh_op_tnl_0')
// (8, 15, 'neigh_op_lft_0')
// (8, 16, 'neigh_op_bnl_0')

wire n363;
// (6, 12, 'sp4_r_v_b_45')
// (6, 13, 'sp4_r_v_b_32')
// (6, 14, 'neigh_op_tnr_4')
// (6, 14, 'sp4_r_v_b_21')
// (6, 15, 'neigh_op_rgt_4')
// (6, 15, 'sp4_r_v_b_8')
// (6, 16, 'neigh_op_bnr_4')
// (7, 11, 'sp4_v_t_45')
// (7, 12, 'sp4_v_b_45')
// (7, 13, 'sp4_v_b_32')
// (7, 14, 'local_g0_4')
// (7, 14, 'local_g0_5')
// (7, 14, 'lutff_1/in_1')
// (7, 14, 'lutff_2/in_0')
// (7, 14, 'lutff_6/in_1')
// (7, 14, 'lutff_7/in_1')
// (7, 14, 'neigh_op_top_4')
// (7, 14, 'sp4_v_b_21')
// (7, 15, 'local_g0_4')
// (7, 15, 'lutff_1/in_1')
// (7, 15, 'lutff_4/out')
// (7, 15, 'lutff_7/in_1')
// (7, 15, 'sp4_v_b_8')
// (7, 16, 'neigh_op_bot_4')
// (8, 14, 'local_g2_4')
// (8, 14, 'local_g3_4')
// (8, 14, 'lutff_0/in_3')
// (8, 14, 'lutff_1/in_2')
// (8, 14, 'lutff_2/in_2')
// (8, 14, 'neigh_op_tnl_4')
// (8, 15, 'neigh_op_lft_4')
// (8, 16, 'neigh_op_bnl_4')

wire n364;
// (6, 13, 'neigh_op_tnr_0')
// (6, 14, 'neigh_op_rgt_0')
// (6, 15, 'neigh_op_bnr_0')
// (7, 11, 'sp4_r_v_b_36')
// (7, 12, 'sp4_r_v_b_25')
// (7, 13, 'local_g0_0')
// (7, 13, 'lutff_6/in_0')
// (7, 13, 'neigh_op_top_0')
// (7, 13, 'sp4_r_v_b_12')
// (7, 14, 'lutff_0/out')
// (7, 14, 'sp4_r_v_b_1')
// (7, 15, 'neigh_op_bot_0')
// (8, 10, 'sp4_v_t_36')
// (8, 11, 'sp4_v_b_36')
// (8, 12, 'local_g2_1')
// (8, 12, 'lutff_3/in_2')
// (8, 12, 'lutff_7/in_2')
// (8, 12, 'sp4_v_b_25')
// (8, 13, 'local_g2_0')
// (8, 13, 'lutff_6/in_0')
// (8, 13, 'neigh_op_tnl_0')
// (8, 13, 'sp4_v_b_12')
// (8, 14, 'neigh_op_lft_0')
// (8, 14, 'sp4_v_b_1')
// (8, 15, 'neigh_op_bnl_0')

wire n365;
// (6, 13, 'neigh_op_tnr_1')
// (6, 14, 'neigh_op_rgt_1')
// (6, 15, 'neigh_op_bnr_1')
// (7, 12, 'sp4_r_v_b_43')
// (7, 13, 'local_g0_1')
// (7, 13, 'local_g0_6')
// (7, 13, 'local_g1_6')
// (7, 13, 'lutff_0/in_3')
// (7, 13, 'lutff_1/in_2')
// (7, 13, 'lutff_3/in_2')
// (7, 13, 'lutff_4/in_2')
// (7, 13, 'neigh_op_top_1')
// (7, 13, 'sp4_r_v_b_30')
// (7, 14, 'lutff_1/out')
// (7, 14, 'sp4_r_v_b_19')
// (7, 15, 'neigh_op_bot_1')
// (7, 15, 'sp4_r_v_b_6')
// (8, 11, 'sp4_v_t_43')
// (8, 12, 'sp4_v_b_43')
// (8, 13, 'neigh_op_tnl_1')
// (8, 13, 'sp4_v_b_30')
// (8, 14, 'neigh_op_lft_1')
// (8, 14, 'sp4_v_b_19')
// (8, 15, 'neigh_op_bnl_1')
// (8, 15, 'sp4_v_b_6')

wire n366;
// (6, 13, 'neigh_op_tnr_2')
// (6, 14, 'neigh_op_rgt_2')
// (6, 15, 'neigh_op_bnr_2')
// (7, 13, 'neigh_op_top_2')
// (7, 14, 'local_g0_2')
// (7, 14, 'local_g1_2')
// (7, 14, 'lutff_0/in_1')
// (7, 14, 'lutff_2/out')
// (7, 14, 'lutff_5/in_1')
// (7, 15, 'neigh_op_bot_2')
// (8, 13, 'neigh_op_tnl_2')
// (8, 14, 'neigh_op_lft_2')
// (8, 15, 'neigh_op_bnl_2')

wire n367;
// (6, 13, 'neigh_op_tnr_4')
// (6, 14, 'neigh_op_rgt_4')
// (6, 15, 'neigh_op_bnr_4')
// (7, 11, 'sp4_r_v_b_44')
// (7, 12, 'local_g2_1')
// (7, 12, 'lutff_1/in_2')
// (7, 12, 'sp4_r_v_b_33')
// (7, 13, 'local_g2_4')
// (7, 13, 'lutff_7/in_3')
// (7, 13, 'neigh_op_top_4')
// (7, 13, 'sp4_r_v_b_20')
// (7, 13, 'sp4_r_v_b_36')
// (7, 14, 'lutff_4/out')
// (7, 14, 'sp4_r_v_b_25')
// (7, 14, 'sp4_r_v_b_9')
// (7, 15, 'neigh_op_bot_4')
// (7, 15, 'sp4_r_v_b_12')
// (7, 16, 'sp4_r_v_b_1')
// (8, 10, 'sp4_v_t_44')
// (8, 11, 'sp4_v_b_44')
// (8, 12, 'sp4_v_b_33')
// (8, 12, 'sp4_v_t_36')
// (8, 13, 'neigh_op_tnl_4')
// (8, 13, 'sp4_v_b_20')
// (8, 13, 'sp4_v_b_36')
// (8, 14, 'neigh_op_lft_4')
// (8, 14, 'sp4_v_b_25')
// (8, 14, 'sp4_v_b_9')
// (8, 15, 'neigh_op_bnl_4')
// (8, 15, 'sp4_v_b_12')
// (8, 16, 'sp4_v_b_1')

wire n368;
// (6, 13, 'neigh_op_tnr_5')
// (6, 14, 'neigh_op_rgt_5')
// (6, 15, 'neigh_op_bnr_5')
// (7, 13, 'local_g1_5')
// (7, 13, 'lutff_6/in_2')
// (7, 13, 'neigh_op_top_5')
// (7, 14, 'lutff_5/out')
// (7, 15, 'neigh_op_bot_5')
// (8, 13, 'neigh_op_tnl_5')
// (8, 14, 'neigh_op_lft_5')
// (8, 15, 'neigh_op_bnl_5')

wire n369;
// (6, 13, 'neigh_op_tnr_6')
// (6, 14, 'neigh_op_rgt_6')
// (6, 15, 'neigh_op_bnr_6')
// (7, 13, 'neigh_op_top_6')
// (7, 14, 'local_g2_6')
// (7, 14, 'local_g3_6')
// (7, 14, 'lutff_3/in_1')
// (7, 14, 'lutff_4/in_1')
// (7, 14, 'lutff_6/out')
// (7, 15, 'neigh_op_bot_6')
// (8, 13, 'neigh_op_tnl_6')
// (8, 14, 'neigh_op_lft_6')
// (8, 15, 'neigh_op_bnl_6')

wire n370;
// (6, 13, 'neigh_op_tnr_7')
// (6, 14, 'neigh_op_rgt_7')
// (6, 15, 'neigh_op_bnr_7')
// (7, 13, 'local_g0_7')
// (7, 13, 'lutff_1/in_0')
// (7, 13, 'lutff_3/in_0')
// (7, 13, 'neigh_op_top_7')
// (7, 14, 'lutff_7/out')
// (7, 15, 'neigh_op_bot_7')
// (8, 13, 'neigh_op_tnl_7')
// (8, 14, 'neigh_op_lft_7')
// (8, 15, 'neigh_op_bnl_7')

reg n371 = 0;
// (6, 13, 'sp4_h_r_11')
// (7, 10, 'sp4_r_v_b_46')
// (7, 11, 'sp4_r_v_b_35')
// (7, 12, 'sp4_r_v_b_22')
// (7, 13, 'sp4_h_r_22')
// (7, 13, 'sp4_r_v_b_11')
// (8, 9, 'sp4_v_t_46')
// (8, 10, 'sp4_v_b_46')
// (8, 11, 'sp4_v_b_35')
// (8, 12, 'local_g0_6')
// (8, 12, 'local_g1_6')
// (8, 12, 'lutff_1/in_3')
// (8, 12, 'lutff_2/in_3')
// (8, 12, 'lutff_4/in_2')
// (8, 12, 'lutff_5/in_1')
// (8, 12, 'lutff_6/in_2')
// (8, 12, 'sp4_v_b_22')
// (8, 13, 'local_g2_3')
// (8, 13, 'lutff_7/in_0')
// (8, 13, 'sp4_h_r_11')
// (8, 13, 'sp4_h_r_35')
// (8, 13, 'sp4_v_b_11')
// (9, 10, 'sp4_r_v_b_38')
// (9, 11, 'sp4_r_v_b_27')
// (9, 12, 'local_g2_6')
// (9, 12, 'lutff_1/in_3')
// (9, 12, 'sp4_r_v_b_14')
// (9, 13, 'local_g1_6')
// (9, 13, 'lutff_2/in_1')
// (9, 13, 'sp4_h_r_22')
// (9, 13, 'sp4_h_r_46')
// (9, 13, 'sp4_r_v_b_3')
// (10, 9, 'sp4_v_t_38')
// (10, 10, 'sp4_v_b_38')
// (10, 11, 'sp4_v_b_27')
// (10, 12, 'neigh_op_tnr_7')
// (10, 12, 'sp4_v_b_14')
// (10, 13, 'neigh_op_rgt_7')
// (10, 13, 'sp4_h_l_46')
// (10, 13, 'sp4_h_r_3')
// (10, 13, 'sp4_h_r_35')
// (10, 13, 'sp4_v_b_3')
// (10, 14, 'neigh_op_bnr_7')
// (11, 12, 'local_g1_7')
// (11, 12, 'lutff_1/in_3')
// (11, 12, 'neigh_op_top_7')
// (11, 13, 'local_g0_7')
// (11, 13, 'lutff_7/in_2')
// (11, 13, 'lutff_7/out')
// (11, 13, 'sp4_h_r_14')
// (11, 13, 'sp4_h_r_46')
// (11, 14, 'neigh_op_bot_7')
// (12, 12, 'neigh_op_tnl_7')
// (12, 13, 'neigh_op_lft_7')
// (12, 13, 'sp4_h_l_46')
// (12, 13, 'sp4_h_r_27')
// (12, 14, 'neigh_op_bnl_7')
// (13, 13, 'span4_horz_27')

wire n372;
// (6, 14, 'neigh_op_tnr_1')
// (6, 15, 'neigh_op_rgt_1')
// (6, 16, 'neigh_op_bnr_1')
// (7, 13, 'sp4_r_v_b_43')
// (7, 14, 'local_g0_6')
// (7, 14, 'local_g1_6')
// (7, 14, 'lutff_4/in_3')
// (7, 14, 'lutff_5/in_3')
// (7, 14, 'neigh_op_top_1')
// (7, 14, 'sp4_r_v_b_30')
// (7, 15, 'lutff_1/out')
// (7, 15, 'sp4_r_v_b_19')
// (7, 16, 'neigh_op_bot_1')
// (7, 16, 'sp4_r_v_b_6')
// (8, 12, 'sp4_v_t_43')
// (8, 13, 'sp4_v_b_43')
// (8, 14, 'neigh_op_tnl_1')
// (8, 14, 'sp4_v_b_30')
// (8, 15, 'neigh_op_lft_1')
// (8, 15, 'sp4_v_b_19')
// (8, 16, 'neigh_op_bnl_1')
// (8, 16, 'sp4_v_b_6')

wire n373;
// (6, 14, 'neigh_op_tnr_2')
// (6, 15, 'neigh_op_rgt_2')
// (6, 16, 'neigh_op_bnr_2')
// (7, 14, 'neigh_op_top_2')
// (7, 15, 'local_g0_2')
// (7, 15, 'lutff_2/out')
// (7, 15, 'lutff_7/in_3')
// (7, 16, 'neigh_op_bot_2')
// (8, 14, 'neigh_op_tnl_2')
// (8, 15, 'neigh_op_lft_2')
// (8, 16, 'neigh_op_bnl_2')

wire n374;
// (6, 14, 'neigh_op_tnr_6')
// (6, 15, 'neigh_op_rgt_6')
// (6, 16, 'neigh_op_bnr_6')
// (7, 14, 'neigh_op_top_6')
// (7, 15, 'local_g1_6')
// (7, 15, 'lutff_1/in_2')
// (7, 15, 'lutff_6/out')
// (7, 15, 'lutff_7/in_2')
// (7, 16, 'neigh_op_bot_6')
// (8, 14, 'neigh_op_tnl_6')
// (8, 15, 'neigh_op_lft_6')
// (8, 16, 'neigh_op_bnl_6')

wire n375;
// (6, 14, 'neigh_op_tnr_7')
// (6, 15, 'neigh_op_rgt_7')
// (6, 16, 'neigh_op_bnr_7')
// (7, 14, 'local_g0_7')
// (7, 14, 'local_g1_7')
// (7, 14, 'lutff_0/in_3')
// (7, 14, 'lutff_3/in_3')
// (7, 14, 'neigh_op_top_7')
// (7, 15, 'lutff_7/out')
// (7, 16, 'neigh_op_bot_7')
// (8, 14, 'neigh_op_tnl_7')
// (8, 15, 'neigh_op_lft_7')
// (8, 16, 'neigh_op_bnl_7')

reg n376 = 0;
// (7, 1, 'sp4_r_v_b_41')
// (7, 2, 'sp4_r_v_b_28')
// (7, 3, 'neigh_op_tnr_2')
// (7, 3, 'sp4_r_v_b_17')
// (7, 4, 'neigh_op_rgt_2')
// (7, 4, 'sp4_r_v_b_4')
// (7, 5, 'neigh_op_bnr_2')
// (8, 0, 'span4_vert_41')
// (8, 1, 'sp4_v_b_41')
// (8, 2, 'sp4_v_b_28')
// (8, 3, 'local_g0_1')
// (8, 3, 'lutff_1/in_0')
// (8, 3, 'lutff_6/in_1')
// (8, 3, 'neigh_op_top_2')
// (8, 3, 'sp4_v_b_17')
// (8, 4, 'lutff_2/out')
// (8, 4, 'sp4_v_b_4')
// (8, 5, 'neigh_op_bot_2')
// (9, 3, 'neigh_op_tnl_2')
// (9, 4, 'neigh_op_lft_2')
// (9, 5, 'neigh_op_bnl_2')

wire n377;
// (7, 2, 'neigh_op_tnr_0')
// (7, 3, 'neigh_op_rgt_0')
// (7, 4, 'neigh_op_bnr_0')
// (7, 4, 'sp4_r_v_b_41')
// (7, 5, 'sp4_r_v_b_28')
// (7, 6, 'sp4_r_v_b_17')
// (7, 7, 'sp4_r_v_b_4')
// (7, 8, 'sp4_r_v_b_42')
// (7, 9, 'local_g0_7')
// (7, 9, 'local_g1_7')
// (7, 9, 'lutff_5/in_2')
// (7, 9, 'lutff_6/in_2')
// (7, 9, 'sp4_r_v_b_31')
// (7, 10, 'sp4_r_v_b_18')
// (7, 11, 'sp4_r_v_b_7')
// (8, 0, 'span12_vert_20')
// (8, 1, 'sp12_v_b_20')
// (8, 2, 'neigh_op_top_0')
// (8, 2, 'sp12_v_b_19')
// (8, 2, 'sp4_r_v_b_44')
// (8, 3, 'lutff_0/out')
// (8, 3, 'sp12_v_b_16')
// (8, 3, 'sp4_r_v_b_33')
// (8, 3, 'sp4_v_t_41')
// (8, 4, 'neigh_op_bot_0')
// (8, 4, 'sp12_v_b_15')
// (8, 4, 'sp4_r_v_b_20')
// (8, 4, 'sp4_v_b_41')
// (8, 5, 'sp12_v_b_12')
// (8, 5, 'sp4_r_v_b_9')
// (8, 5, 'sp4_v_b_28')
// (8, 6, 'sp12_v_b_11')
// (8, 6, 'sp4_r_v_b_44')
// (8, 6, 'sp4_v_b_17')
// (8, 7, 'sp12_v_b_8')
// (8, 7, 'sp4_r_v_b_33')
// (8, 7, 'sp4_v_b_4')
// (8, 7, 'sp4_v_t_42')
// (8, 8, 'sp12_v_b_7')
// (8, 8, 'sp4_r_v_b_20')
// (8, 8, 'sp4_v_b_42')
// (8, 9, 'local_g3_4')
// (8, 9, 'lutff_0/in_1')
// (8, 9, 'lutff_1/in_2')
// (8, 9, 'sp12_v_b_4')
// (8, 9, 'sp4_r_v_b_9')
// (8, 9, 'sp4_v_b_31')
// (8, 10, 'sp12_v_b_3')
// (8, 10, 'sp4_v_b_18')
// (8, 11, 'sp12_v_b_0')
// (8, 11, 'sp4_v_b_7')
// (9, 1, 'sp4_v_t_44')
// (9, 2, 'neigh_op_tnl_0')
// (9, 2, 'sp4_v_b_44')
// (9, 3, 'neigh_op_lft_0')
// (9, 3, 'sp4_v_b_33')
// (9, 4, 'neigh_op_bnl_0')
// (9, 4, 'sp4_v_b_20')
// (9, 5, 'sp4_v_b_9')
// (9, 5, 'sp4_v_t_44')
// (9, 6, 'sp4_v_b_44')
// (9, 7, 'sp4_v_b_33')
// (9, 8, 'sp4_v_b_20')
// (9, 9, 'local_g0_1')
// (9, 9, 'lutff_5/in_2')
// (9, 9, 'sp4_v_b_9')

wire n378;
// (7, 2, 'neigh_op_tnr_1')
// (7, 3, 'neigh_op_rgt_1')
// (7, 4, 'neigh_op_bnr_1')
// (8, 2, 'neigh_op_top_1')
// (8, 3, 'local_g2_1')
// (8, 3, 'lutff_0/in_3')
// (8, 3, 'lutff_1/out')
// (8, 4, 'neigh_op_bot_1')
// (9, 2, 'neigh_op_tnl_1')
// (9, 3, 'neigh_op_lft_1')
// (9, 4, 'neigh_op_bnl_1')

reg n379 = 0;
// (7, 2, 'neigh_op_tnr_2')
// (7, 3, 'neigh_op_rgt_2')
// (7, 4, 'neigh_op_bnr_2')
// (8, 2, 'neigh_op_top_2')
// (8, 3, 'local_g1_2')
// (8, 3, 'lutff_0/in_1')
// (8, 3, 'lutff_2/out')
// (8, 4, 'neigh_op_bot_2')
// (9, 2, 'neigh_op_tnl_2')
// (9, 3, 'local_g1_2')
// (9, 3, 'lutff_4/in_1')
// (9, 3, 'neigh_op_lft_2')
// (9, 4, 'neigh_op_bnl_2')

reg n380 = 0;
// (7, 2, 'neigh_op_tnr_3')
// (7, 3, 'neigh_op_rgt_3')
// (7, 4, 'neigh_op_bnr_3')
// (8, 2, 'neigh_op_top_3')
// (8, 3, 'lutff_3/out')
// (8, 4, 'local_g1_3')
// (8, 4, 'lutff_4/in_0')
// (8, 4, 'neigh_op_bot_3')
// (9, 2, 'neigh_op_tnl_3')
// (9, 3, 'neigh_op_lft_3')
// (9, 4, 'neigh_op_bnl_3')

reg n381 = 0;
// (7, 2, 'neigh_op_tnr_4')
// (7, 3, 'neigh_op_rgt_4')
// (7, 4, 'neigh_op_bnr_4')
// (8, 2, 'neigh_op_top_4')
// (8, 3, 'local_g1_4')
// (8, 3, 'lutff_4/out')
// (8, 3, 'lutff_7/in_0')
// (8, 4, 'neigh_op_bot_4')
// (9, 2, 'neigh_op_tnl_4')
// (9, 3, 'neigh_op_lft_4')
// (9, 4, 'neigh_op_bnl_4')

reg n382 = 0;
// (7, 2, 'neigh_op_tnr_6')
// (7, 3, 'neigh_op_rgt_6')
// (7, 4, 'neigh_op_bnr_6')
// (8, 2, 'neigh_op_top_6')
// (8, 3, 'local_g0_6')
// (8, 3, 'lutff_4/in_0')
// (8, 3, 'lutff_6/out')
// (8, 4, 'neigh_op_bot_6')
// (9, 2, 'neigh_op_tnl_6')
// (9, 3, 'neigh_op_lft_6')
// (9, 4, 'neigh_op_bnl_6')

reg n383 = 0;
// (7, 2, 'neigh_op_tnr_7')
// (7, 3, 'neigh_op_rgt_7')
// (7, 4, 'neigh_op_bnr_7')
// (8, 2, 'neigh_op_top_7')
// (8, 3, 'local_g1_7')
// (8, 3, 'lutff_2/in_0')
// (8, 3, 'lutff_7/out')
// (8, 4, 'neigh_op_bot_7')
// (9, 2, 'neigh_op_tnl_7')
// (9, 3, 'neigh_op_lft_7')
// (9, 4, 'neigh_op_bnl_7')

reg n384 = 0;
// (7, 2, 'sp4_r_v_b_38')
// (7, 3, 'neigh_op_tnr_7')
// (7, 3, 'sp4_r_v_b_27')
// (7, 3, 'sp4_r_v_b_43')
// (7, 4, 'neigh_op_rgt_7')
// (7, 4, 'sp4_r_v_b_14')
// (7, 4, 'sp4_r_v_b_30')
// (7, 5, 'neigh_op_bnr_7')
// (7, 5, 'sp4_r_v_b_19')
// (7, 5, 'sp4_r_v_b_3')
// (7, 6, 'sp4_r_v_b_6')
// (8, 1, 'sp4_v_t_38')
// (8, 2, 'sp4_v_b_38')
// (8, 2, 'sp4_v_t_43')
// (8, 3, 'neigh_op_top_7')
// (8, 3, 'sp4_v_b_27')
// (8, 3, 'sp4_v_b_43')
// (8, 4, 'lutff_7/out')
// (8, 4, 'sp4_v_b_14')
// (8, 4, 'sp4_v_b_30')
// (8, 5, 'local_g1_3')
// (8, 5, 'lutff_5/in_1')
// (8, 5, 'neigh_op_bot_7')
// (8, 5, 'sp4_v_b_19')
// (8, 5, 'sp4_v_b_3')
// (8, 6, 'local_g1_6')
// (8, 6, 'lutff_2/in_1')
// (8, 6, 'sp4_v_b_6')
// (9, 3, 'neigh_op_tnl_7')
// (9, 4, 'neigh_op_lft_7')
// (9, 5, 'neigh_op_bnl_7')

reg n385 = 0;
// (7, 3, 'neigh_op_tnr_0')
// (7, 4, 'neigh_op_rgt_0')
// (7, 5, 'neigh_op_bnr_0')
// (8, 3, 'neigh_op_top_0')
// (8, 4, 'local_g1_0')
// (8, 4, 'lutff_0/out')
// (8, 4, 'lutff_7/in_0')
// (8, 5, 'neigh_op_bot_0')
// (9, 3, 'neigh_op_tnl_0')
// (9, 4, 'neigh_op_lft_0')
// (9, 5, 'neigh_op_bnl_0')

reg n386 = 0;
// (7, 3, 'neigh_op_tnr_4')
// (7, 4, 'neigh_op_rgt_4')
// (7, 5, 'neigh_op_bnr_4')
// (8, 3, 'neigh_op_top_4')
// (8, 4, 'local_g1_4')
// (8, 4, 'lutff_4/out')
// (8, 4, 'lutff_5/in_0')
// (8, 5, 'neigh_op_bot_4')
// (9, 3, 'neigh_op_tnl_4')
// (9, 4, 'neigh_op_lft_4')
// (9, 5, 'neigh_op_bnl_4')

reg n387 = 0;
// (7, 3, 'neigh_op_tnr_5')
// (7, 4, 'neigh_op_rgt_5')
// (7, 5, 'neigh_op_bnr_5')
// (8, 3, 'neigh_op_top_5')
// (8, 4, 'local_g1_5')
// (8, 4, 'lutff_2/in_0')
// (8, 4, 'lutff_5/out')
// (8, 5, 'neigh_op_bot_5')
// (9, 3, 'neigh_op_tnl_5')
// (9, 4, 'neigh_op_lft_5')
// (9, 5, 'neigh_op_bnl_5')

reg n388 = 0;
// (7, 4, 'neigh_op_tnr_0')
// (7, 5, 'neigh_op_rgt_0')
// (7, 6, 'neigh_op_bnr_0')
// (8, 4, 'local_g0_0')
// (8, 4, 'lutff_0/in_0')
// (8, 4, 'neigh_op_top_0')
// (8, 5, 'lutff_0/out')
// (8, 6, 'neigh_op_bot_0')
// (9, 4, 'neigh_op_tnl_0')
// (9, 5, 'neigh_op_lft_0')
// (9, 6, 'neigh_op_bnl_0')

reg n389 = 0;
// (7, 4, 'neigh_op_tnr_1')
// (7, 5, 'neigh_op_rgt_1')
// (7, 6, 'neigh_op_bnr_1')
// (8, 4, 'neigh_op_top_1')
// (8, 5, 'local_g0_1')
// (8, 5, 'lutff_1/out')
// (8, 5, 'lutff_3/in_0')
// (8, 6, 'neigh_op_bot_1')
// (9, 4, 'neigh_op_tnl_1')
// (9, 5, 'neigh_op_lft_1')
// (9, 6, 'neigh_op_bnl_1')

reg n390 = 0;
// (7, 4, 'neigh_op_tnr_2')
// (7, 5, 'neigh_op_rgt_2')
// (7, 6, 'neigh_op_bnr_2')
// (8, 4, 'neigh_op_top_2')
// (8, 5, 'local_g0_2')
// (8, 5, 'lutff_2/out')
// (8, 5, 'lutff_4/in_0')
// (8, 6, 'neigh_op_bot_2')
// (9, 4, 'neigh_op_tnl_2')
// (9, 5, 'neigh_op_lft_2')
// (9, 6, 'neigh_op_bnl_2')

reg n391 = 0;
// (7, 4, 'neigh_op_tnr_3')
// (7, 5, 'neigh_op_rgt_3')
// (7, 6, 'neigh_op_bnr_3')
// (8, 4, 'neigh_op_top_3')
// (8, 5, 'local_g0_3')
// (8, 5, 'lutff_3/out')
// (8, 5, 'lutff_6/in_1')
// (8, 6, 'local_g0_3')
// (8, 6, 'lutff_1/in_0')
// (8, 6, 'neigh_op_bot_3')
// (9, 4, 'neigh_op_tnl_3')
// (9, 5, 'neigh_op_lft_3')
// (9, 6, 'neigh_op_bnl_3')

reg n392 = 0;
// (7, 4, 'neigh_op_tnr_4')
// (7, 5, 'neigh_op_rgt_4')
// (7, 6, 'neigh_op_bnr_4')
// (8, 4, 'neigh_op_top_4')
// (8, 5, 'local_g0_4')
// (8, 5, 'local_g1_4')
// (8, 5, 'lutff_4/out')
// (8, 5, 'lutff_5/in_0')
// (8, 5, 'lutff_6/in_0')
// (8, 6, 'local_g0_4')
// (8, 6, 'lutff_1/in_1')
// (8, 6, 'lutff_4/in_2')
// (8, 6, 'neigh_op_bot_4')
// (9, 4, 'neigh_op_tnl_4')
// (9, 5, 'neigh_op_lft_4')
// (9, 6, 'neigh_op_bnl_4')

reg n393 = 0;
// (7, 4, 'neigh_op_tnr_5')
// (7, 5, 'neigh_op_rgt_5')
// (7, 6, 'neigh_op_bnr_5')
// (8, 4, 'neigh_op_top_5')
// (8, 5, 'local_g0_5')
// (8, 5, 'lutff_5/out')
// (8, 5, 'lutff_7/in_0')
// (8, 6, 'neigh_op_bot_5')
// (9, 4, 'neigh_op_tnl_5')
// (9, 5, 'neigh_op_lft_5')
// (9, 6, 'neigh_op_bnl_5')

reg n394 = 0;
// (7, 4, 'neigh_op_tnr_6')
// (7, 5, 'neigh_op_rgt_6')
// (7, 6, 'neigh_op_bnr_6')
// (8, 4, 'neigh_op_top_6')
// (8, 5, 'local_g0_6')
// (8, 5, 'lutff_0/in_0')
// (8, 5, 'lutff_6/out')
// (8, 6, 'neigh_op_bot_6')
// (9, 4, 'neigh_op_tnl_6')
// (9, 5, 'neigh_op_lft_6')
// (9, 6, 'neigh_op_bnl_6')

reg n395 = 0;
// (7, 4, 'neigh_op_tnr_7')
// (7, 5, 'neigh_op_rgt_7')
// (7, 6, 'neigh_op_bnr_7')
// (8, 4, 'neigh_op_top_7')
// (8, 5, 'local_g1_7')
// (8, 5, 'lutff_2/in_0')
// (8, 5, 'lutff_7/out')
// (8, 6, 'neigh_op_bot_7')
// (9, 4, 'neigh_op_tnl_7')
// (9, 5, 'neigh_op_lft_7')
// (9, 6, 'neigh_op_bnl_7')

wire n396;
// (7, 5, 'neigh_op_tnr_1')
// (7, 6, 'neigh_op_rgt_1')
// (7, 7, 'neigh_op_bnr_1')
// (8, 5, 'neigh_op_top_1')
// (8, 6, 'local_g2_1')
// (8, 6, 'lutff_1/out')
// (8, 6, 'lutff_2/in_3')
// (8, 7, 'neigh_op_bot_1')
// (9, 5, 'neigh_op_tnl_1')
// (9, 6, 'neigh_op_lft_1')
// (9, 7, 'neigh_op_bnl_1')

wire n397;
// (7, 5, 'neigh_op_tnr_2')
// (7, 6, 'neigh_op_rgt_2')
// (7, 7, 'neigh_op_bnr_2')
// (8, 4, 'sp12_v_t_23')
// (8, 4, 'sp4_r_v_b_45')
// (8, 5, 'neigh_op_top_2')
// (8, 5, 'sp12_v_b_23')
// (8, 5, 'sp4_r_v_b_32')
// (8, 6, 'lutff_2/out')
// (8, 6, 'sp12_v_b_20')
// (8, 6, 'sp4_r_v_b_21')
// (8, 7, 'neigh_op_bot_2')
// (8, 7, 'sp12_v_b_19')
// (8, 7, 'sp4_r_v_b_8')
// (8, 8, 'sp12_v_b_16')
// (8, 8, 'sp4_r_v_b_45')
// (8, 9, 'local_g2_7')
// (8, 9, 'lutff_0/in_3')
// (8, 9, 'sp12_v_b_15')
// (8, 9, 'sp4_r_v_b_32')
// (8, 10, 'local_g2_4')
// (8, 10, 'lutff_7/in_3')
// (8, 10, 'sp12_v_b_12')
// (8, 10, 'sp4_r_v_b_21')
// (8, 11, 'sp12_v_b_11')
// (8, 11, 'sp4_r_v_b_8')
// (8, 12, 'sp12_v_b_8')
// (8, 13, 'sp12_v_b_7')
// (8, 14, 'sp12_v_b_4')
// (8, 15, 'sp12_v_b_3')
// (8, 16, 'sp12_v_b_0')
// (9, 3, 'sp4_v_t_45')
// (9, 4, 'sp4_v_b_45')
// (9, 5, 'neigh_op_tnl_2')
// (9, 5, 'sp4_v_b_32')
// (9, 6, 'neigh_op_lft_2')
// (9, 6, 'sp4_v_b_21')
// (9, 7, 'local_g1_0')
// (9, 7, 'lutff_0/in_3')
// (9, 7, 'neigh_op_bnl_2')
// (9, 7, 'sp4_v_b_8')
// (9, 7, 'sp4_v_t_45')
// (9, 8, 'sp4_v_b_45')
// (9, 9, 'local_g2_0')
// (9, 9, 'lutff_0/in_2')
// (9, 9, 'sp4_v_b_32')
// (9, 10, 'local_g1_5')
// (9, 10, 'lutff_0/in_2')
// (9, 10, 'sp4_v_b_21')
// (9, 11, 'sp4_v_b_8')

reg n398 = 0;
// (7, 5, 'neigh_op_tnr_4')
// (7, 6, 'neigh_op_rgt_4')
// (7, 7, 'neigh_op_bnr_4')
// (8, 5, 'neigh_op_top_4')
// (8, 6, 'local_g1_4')
// (8, 6, 'lutff_4/out')
// (8, 6, 'lutff_7/in_0')
// (8, 7, 'neigh_op_bot_4')
// (9, 5, 'neigh_op_tnl_4')
// (9, 6, 'neigh_op_lft_4')
// (9, 7, 'neigh_op_bnl_4')

reg \d_out[0] = 0 ;
// (7, 5, 'neigh_op_tnr_5')
// (7, 6, 'neigh_op_rgt_5')
// (7, 7, 'neigh_op_bnr_5')
// (8, 1, 'sp4_r_v_b_43')
// (8, 2, 'sp4_r_v_b_30')
// (8, 3, 'sp4_r_v_b_19')
// (8, 4, 'sp4_r_v_b_6')
// (8, 5, 'neigh_op_top_5')
// (8, 5, 'sp4_r_v_b_38')
// (8, 6, 'lutff_5/out')
// (8, 6, 'sp4_r_v_b_27')
// (8, 7, 'neigh_op_bot_5')
// (8, 7, 'sp4_r_v_b_14')
// (8, 8, 'sp4_r_v_b_3')
// (9, 0, 'io_1/D_OUT_0')
// (9, 0, 'io_1/PAD')
// (9, 0, 'local_g0_3')
// (9, 0, 'span4_vert_43')
// (9, 1, 'sp4_v_b_43')
// (9, 2, 'sp4_v_b_30')
// (9, 3, 'sp4_v_b_19')
// (9, 4, 'sp4_v_b_6')
// (9, 4, 'sp4_v_t_38')
// (9, 5, 'neigh_op_tnl_5')
// (9, 5, 'sp4_v_b_38')
// (9, 6, 'neigh_op_lft_5')
// (9, 6, 'sp4_v_b_27')
// (9, 7, 'neigh_op_bnl_5')
// (9, 7, 'sp4_v_b_14')
// (9, 8, 'sp4_v_b_3')

reg n400 = 0;
// (7, 5, 'neigh_op_tnr_6')
// (7, 6, 'neigh_op_rgt_6')
// (7, 7, 'neigh_op_bnr_6')
// (8, 5, 'neigh_op_top_6')
// (8, 6, 'lutff_6/out')
// (8, 7, 'local_g0_6')
// (8, 7, 'lutff_6/in_0')
// (8, 7, 'neigh_op_bot_6')
// (9, 5, 'neigh_op_tnl_6')
// (9, 6, 'neigh_op_lft_6')
// (9, 7, 'neigh_op_bnl_6')

reg n401 = 0;
// (7, 5, 'neigh_op_tnr_7')
// (7, 6, 'neigh_op_rgt_7')
// (7, 7, 'neigh_op_bnr_7')
// (8, 5, 'local_g0_7')
// (8, 5, 'lutff_1/in_0')
// (8, 5, 'neigh_op_top_7')
// (8, 6, 'lutff_7/out')
// (8, 7, 'neigh_op_bot_7')
// (9, 5, 'neigh_op_tnl_7')
// (9, 6, 'neigh_op_lft_7')
// (9, 7, 'neigh_op_bnl_7')

wire n402;
// (7, 6, 'neigh_op_tnr_0')
// (7, 7, 'neigh_op_rgt_0')
// (7, 8, 'neigh_op_bnr_0')
// (8, 6, 'neigh_op_top_0')
// (8, 7, 'lutff_0/out')
// (8, 8, 'neigh_op_bot_0')
// (9, 6, 'local_g2_0')
// (9, 6, 'local_g3_0')
// (9, 6, 'lutff_0/in_0')
// (9, 6, 'lutff_4/in_1')
// (9, 6, 'neigh_op_tnl_0')
// (9, 7, 'neigh_op_lft_0')
// (9, 8, 'neigh_op_bnl_0')

reg n403 = 0;
// (7, 6, 'neigh_op_tnr_1')
// (7, 7, 'neigh_op_rgt_1')
// (7, 8, 'neigh_op_bnr_1')
// (8, 0, 'span12_vert_14')
// (8, 1, 'sp12_v_b_14')
// (8, 2, 'sp12_v_b_13')
// (8, 3, 'sp12_v_b_10')
// (8, 4, 'sp12_v_b_9')
// (8, 5, 'sp12_v_b_6')
// (8, 6, 'neigh_op_top_1')
// (8, 6, 'sp12_v_b_5')
// (8, 7, 'local_g1_1')
// (8, 7, 'lutff_1/out')
// (8, 7, 'lutff_3/in_1')
// (8, 7, 'sp12_v_b_2')
// (8, 8, 'neigh_op_bot_1')
// (8, 8, 'sp12_h_r_1')
// (8, 8, 'sp12_v_b_1')
// (9, 6, 'neigh_op_tnl_1')
// (9, 7, 'neigh_op_lft_1')
// (9, 8, 'neigh_op_bnl_1')
// (9, 8, 'sp12_h_r_2')
// (10, 8, 'sp12_h_r_5')
// (11, 8, 'local_g1_6')
// (11, 8, 'lutff_3/in_0')
// (11, 8, 'sp12_h_r_6')
// (12, 8, 'sp12_h_r_9')
// (13, 8, 'span12_horz_9')

reg n404 = 0;
// (7, 6, 'neigh_op_tnr_6')
// (7, 7, 'neigh_op_rgt_6')
// (7, 8, 'neigh_op_bnr_6')
// (8, 6, 'neigh_op_top_6')
// (8, 7, 'lutff_6/out')
// (8, 8, 'local_g1_6')
// (8, 8, 'lutff_3/in_0')
// (8, 8, 'neigh_op_bot_6')
// (9, 6, 'neigh_op_tnl_6')
// (9, 7, 'neigh_op_lft_6')
// (9, 8, 'neigh_op_bnl_6')

reg n405 = 0;
// (7, 6, 'neigh_op_tnr_7')
// (7, 7, 'neigh_op_rgt_7')
// (7, 8, 'neigh_op_bnr_7')
// (8, 6, 'neigh_op_top_7')
// (8, 7, 'local_g1_7')
// (8, 7, 'lutff_0/in_0')
// (8, 7, 'lutff_1/in_1')
// (8, 7, 'lutff_7/out')
// (8, 8, 'neigh_op_bot_7')
// (9, 6, 'neigh_op_tnl_7')
// (9, 7, 'neigh_op_lft_7')
// (9, 8, 'neigh_op_bnl_7')

wire n406;
// (7, 6, 'sp4_r_v_b_40')
// (7, 7, 'neigh_op_tnr_0')
// (7, 7, 'sp4_r_v_b_29')
// (7, 8, 'neigh_op_rgt_0')
// (7, 8, 'sp4_r_v_b_16')
// (7, 9, 'neigh_op_bnr_0')
// (7, 9, 'sp4_r_v_b_5')
// (8, 5, 'sp4_v_t_40')
// (8, 6, 'sp4_v_b_40')
// (8, 7, 'neigh_op_top_0')
// (8, 7, 'sp4_v_b_29')
// (8, 8, 'local_g0_0')
// (8, 8, 'lutff_0/out')
// (8, 8, 'lutff_4/in_2')
// (8, 8, 'sp4_h_r_0')
// (8, 8, 'sp4_v_b_16')
// (8, 9, 'neigh_op_bot_0')
// (8, 9, 'sp4_h_r_5')
// (8, 9, 'sp4_v_b_5')
// (9, 7, 'neigh_op_tnl_0')
// (9, 8, 'neigh_op_lft_0')
// (9, 8, 'sp4_h_r_13')
// (9, 9, 'neigh_op_bnl_0')
// (9, 9, 'sp4_h_r_16')
// (10, 8, 'sp4_h_r_24')
// (10, 9, 'sp4_h_r_29')
// (11, 8, 'sp4_h_r_37')
// (11, 9, 'local_g2_0')
// (11, 9, 'local_g2_5')
// (11, 9, 'lutff_4/in_3')
// (11, 9, 'lutff_5/in_3')
// (11, 9, 'lutff_6/in_3')
// (11, 9, 'sp4_h_r_40')
// (11, 9, 'sp4_r_v_b_37')
// (11, 10, 'sp4_r_v_b_24')
// (11, 11, 'sp4_r_v_b_13')
// (11, 12, 'sp4_r_v_b_0')
// (12, 8, 'sp4_h_l_37')
// (12, 8, 'sp4_v_t_37')
// (12, 9, 'sp4_h_l_40')
// (12, 9, 'sp4_v_b_37')
// (12, 10, 'sp4_v_b_24')
// (12, 11, 'sp4_v_b_13')
// (12, 12, 'sp4_v_b_0')

wire n407;
// (7, 6, 'sp4_r_v_b_47')
// (7, 7, 'sp4_r_v_b_34')
// (7, 8, 'neigh_op_tnr_5')
// (7, 8, 'sp4_r_v_b_23')
// (7, 9, 'neigh_op_rgt_5')
// (7, 9, 'sp4_r_v_b_10')
// (7, 10, 'neigh_op_bnr_5')
// (8, 5, 'sp4_v_t_47')
// (8, 6, 'sp4_v_b_47')
// (8, 7, 'local_g2_2')
// (8, 7, 'lutff_1/in_3')
// (8, 7, 'lutff_3/in_3')
// (8, 7, 'sp4_v_b_34')
// (8, 8, 'local_g1_5')
// (8, 8, 'lutff_0/in_2')
// (8, 8, 'neigh_op_top_5')
// (8, 8, 'sp4_v_b_23')
// (8, 9, 'lutff_5/out')
// (8, 9, 'sp4_v_b_10')
// (8, 10, 'neigh_op_bot_5')
// (9, 8, 'neigh_op_tnl_5')
// (9, 9, 'neigh_op_lft_5')
// (9, 10, 'neigh_op_bnl_5')

reg n408 = 0;
// (7, 7, 'neigh_op_tnr_1')
// (7, 8, 'neigh_op_rgt_1')
// (7, 9, 'neigh_op_bnr_1')
// (8, 7, 'neigh_op_top_1')
// (8, 8, 'local_g2_1')
// (8, 8, 'lutff_1/out')
// (8, 8, 'lutff_7/in_0')
// (8, 9, 'neigh_op_bot_1')
// (9, 7, 'neigh_op_tnl_1')
// (9, 8, 'neigh_op_lft_1')
// (9, 9, 'neigh_op_bnl_1')

reg n409 = 0;
// (7, 7, 'neigh_op_tnr_2')
// (7, 8, 'neigh_op_rgt_2')
// (7, 9, 'local_g0_2')
// (7, 9, 'lutff_7/in_3')
// (7, 9, 'neigh_op_bnr_2')
// (8, 7, 'neigh_op_top_2')
// (8, 8, 'local_g0_2')
// (8, 8, 'local_g1_2')
// (8, 8, 'lutff_2/out')
// (8, 8, 'lutff_4/in_3')
// (8, 8, 'lutff_6/in_2')
// (8, 9, 'neigh_op_bot_2')
// (9, 7, 'neigh_op_tnl_2')
// (9, 8, 'neigh_op_lft_2')
// (9, 9, 'neigh_op_bnl_2')

reg n410 = 0;
// (7, 7, 'neigh_op_tnr_3')
// (7, 8, 'neigh_op_rgt_3')
// (7, 9, 'neigh_op_bnr_3')
// (8, 7, 'neigh_op_top_3')
// (8, 8, 'local_g0_3')
// (8, 8, 'lutff_3/out')
// (8, 8, 'lutff_5/in_0')
// (8, 9, 'neigh_op_bot_3')
// (9, 7, 'neigh_op_tnl_3')
// (9, 8, 'neigh_op_lft_3')
// (9, 9, 'neigh_op_bnl_3')

reg \d_out[2] = 0 ;
// (7, 7, 'neigh_op_tnr_4')
// (7, 8, 'neigh_op_rgt_4')
// (7, 9, 'neigh_op_bnr_4')
// (8, 0, 'io_1/D_OUT_0')
// (8, 0, 'io_1/PAD')
// (8, 0, 'local_g0_7')
// (8, 0, 'span12_vert_23')
// (8, 1, 'sp12_v_b_23')
// (8, 2, 'sp12_v_b_20')
// (8, 3, 'sp12_v_b_19')
// (8, 4, 'sp12_v_b_16')
// (8, 5, 'sp12_v_b_15')
// (8, 6, 'sp12_v_b_12')
// (8, 7, 'neigh_op_top_4')
// (8, 7, 'sp12_v_b_11')
// (8, 8, 'lutff_4/out')
// (8, 8, 'sp12_v_b_8')
// (8, 9, 'neigh_op_bot_4')
// (8, 9, 'sp12_v_b_7')
// (8, 10, 'sp12_v_b_4')
// (8, 11, 'sp12_v_b_3')
// (8, 12, 'sp12_v_b_0')
// (9, 7, 'neigh_op_tnl_4')
// (9, 8, 'neigh_op_lft_4')
// (9, 9, 'neigh_op_bnl_4')

reg n412 = 0;
// (7, 7, 'neigh_op_tnr_5')
// (7, 8, 'neigh_op_rgt_5')
// (7, 9, 'neigh_op_bnr_5')
// (8, 1, 'sp12_v_t_22')
// (8, 2, 'sp12_v_b_22')
// (8, 3, 'sp12_v_b_21')
// (8, 4, 'sp12_v_b_18')
// (8, 5, 'sp12_v_b_17')
// (8, 6, 'sp12_v_b_14')
// (8, 7, 'neigh_op_top_5')
// (8, 7, 'sp12_v_b_13')
// (8, 8, 'lutff_5/out')
// (8, 8, 'sp12_v_b_10')
// (8, 9, 'neigh_op_bot_5')
// (8, 9, 'sp12_v_b_9')
// (8, 10, 'sp12_v_b_6')
// (8, 11, 'sp12_v_b_5')
// (8, 12, 'local_g3_2')
// (8, 12, 'lutff_0/in_3')
// (8, 12, 'sp12_v_b_2')
// (8, 13, 'sp12_v_b_1')
// (9, 7, 'neigh_op_tnl_5')
// (9, 8, 'neigh_op_lft_5')
// (9, 9, 'neigh_op_bnl_5')

reg n413 = 0;
// (7, 7, 'neigh_op_tnr_6')
// (7, 8, 'neigh_op_rgt_6')
// (7, 9, 'neigh_op_bnr_6')
// (8, 7, 'neigh_op_top_6')
// (8, 8, 'local_g3_6')
// (8, 8, 'lutff_1/in_0')
// (8, 8, 'lutff_6/out')
// (8, 9, 'neigh_op_bot_6')
// (9, 7, 'neigh_op_tnl_6')
// (9, 8, 'neigh_op_lft_6')
// (9, 9, 'neigh_op_bnl_6')

reg n414 = 0;
// (7, 7, 'neigh_op_tnr_7')
// (7, 8, 'neigh_op_rgt_7')
// (7, 9, 'neigh_op_bnr_7')
// (8, 7, 'neigh_op_top_7')
// (8, 8, 'local_g1_7')
// (8, 8, 'lutff_2/in_0')
// (8, 8, 'lutff_7/out')
// (8, 9, 'neigh_op_bot_7')
// (9, 7, 'neigh_op_tnl_7')
// (9, 8, 'neigh_op_lft_7')
// (9, 9, 'neigh_op_bnl_7')

wire n415;
// (7, 7, 'sp4_r_v_b_40')
// (7, 8, 'neigh_op_tnr_0')
// (7, 8, 'sp4_r_v_b_29')
// (7, 9, 'neigh_op_rgt_0')
// (7, 9, 'sp4_r_v_b_16')
// (7, 10, 'neigh_op_bnr_0')
// (7, 10, 'sp4_r_v_b_5')
// (8, 6, 'sp4_v_t_40')
// (8, 7, 'sp4_v_b_40')
// (8, 8, 'neigh_op_top_0')
// (8, 8, 'sp4_v_b_29')
// (8, 9, 'lutff_0/out')
// (8, 9, 'sp4_v_b_16')
// (8, 10, 'local_g0_0')
// (8, 10, 'local_g0_5')
// (8, 10, 'local_g1_3')
// (8, 10, 'lutff_0/in_1')
// (8, 10, 'lutff_1/in_3')
// (8, 10, 'lutff_2/in_3')
// (8, 10, 'lutff_5/in_1')
// (8, 10, 'neigh_op_bot_0')
// (8, 10, 'sp4_h_r_11')
// (8, 10, 'sp4_v_b_5')
// (9, 8, 'neigh_op_tnl_0')
// (9, 9, 'neigh_op_lft_0')
// (9, 10, 'neigh_op_bnl_0')
// (9, 10, 'sp4_h_r_22')
// (10, 10, 'sp4_h_r_35')
// (11, 10, 'sp4_h_r_46')
// (12, 10, 'sp4_h_l_46')

wire n416;
// (7, 8, 'neigh_op_tnr_1')
// (7, 9, 'neigh_op_rgt_1')
// (7, 10, 'neigh_op_bnr_1')
// (8, 6, 'sp12_v_t_22')
// (8, 6, 'sp4_r_v_b_38')
// (8, 7, 'sp12_v_b_22')
// (8, 7, 'sp4_r_v_b_27')
// (8, 7, 'sp4_r_v_b_43')
// (8, 8, 'neigh_op_top_1')
// (8, 8, 'sp12_v_b_21')
// (8, 8, 'sp4_r_v_b_14')
// (8, 8, 'sp4_r_v_b_30')
// (8, 9, 'lutff_1/out')
// (8, 9, 'sp12_v_b_18')
// (8, 9, 'sp4_r_v_b_19')
// (8, 9, 'sp4_r_v_b_3')
// (8, 10, 'local_g0_1')
// (8, 10, 'lutff_4/in_1')
// (8, 10, 'lutff_7/in_2')
// (8, 10, 'neigh_op_bot_1')
// (8, 10, 'sp12_v_b_17')
// (8, 10, 'sp4_r_v_b_6')
// (8, 11, 'local_g2_6')
// (8, 11, 'lutff_5/in_3')
// (8, 11, 'sp12_v_b_14')
// (8, 11, 'sp4_r_v_b_44')
// (8, 12, 'sp12_v_b_13')
// (8, 12, 'sp4_r_v_b_33')
// (8, 13, 'sp12_v_b_10')
// (8, 13, 'sp4_r_v_b_20')
// (8, 14, 'sp12_v_b_9')
// (8, 14, 'sp4_r_v_b_9')
// (8, 15, 'sp12_v_b_6')
// (8, 16, 'sp12_v_b_5')
// (8, 17, 'span12_vert_2')
// (9, 5, 'sp4_v_t_38')
// (9, 6, 'sp4_v_b_38')
// (9, 6, 'sp4_v_t_43')
// (9, 7, 'sp4_v_b_27')
// (9, 7, 'sp4_v_b_43')
// (9, 8, 'neigh_op_tnl_1')
// (9, 8, 'sp4_v_b_14')
// (9, 8, 'sp4_v_b_30')
// (9, 9, 'local_g0_3')
// (9, 9, 'lutff_4/in_1')
// (9, 9, 'neigh_op_lft_1')
// (9, 9, 'sp4_v_b_19')
// (9, 9, 'sp4_v_b_3')
// (9, 10, 'local_g1_6')
// (9, 10, 'lutff_0/in_3')
// (9, 10, 'neigh_op_bnl_1')
// (9, 10, 'sp4_v_b_6')
// (9, 10, 'sp4_v_t_44')
// (9, 11, 'local_g2_4')
// (9, 11, 'local_g3_4')
// (9, 11, 'lutff_0/in_2')
// (9, 11, 'lutff_3/in_2')
// (9, 11, 'sp4_v_b_44')
// (9, 12, 'sp4_v_b_33')
// (9, 13, 'sp4_v_b_20')
// (9, 14, 'sp4_v_b_9')

wire n417;
// (7, 8, 'neigh_op_tnr_4')
// (7, 9, 'neigh_op_rgt_4')
// (7, 10, 'neigh_op_bnr_4')
// (8, 8, 'neigh_op_top_4')
// (8, 9, 'local_g1_4')
// (8, 9, 'lutff_4/out')
// (8, 9, 'lutff_7/in_0')
// (8, 10, 'neigh_op_bot_4')
// (9, 8, 'neigh_op_tnl_4')
// (9, 9, 'neigh_op_lft_4')
// (9, 10, 'neigh_op_bnl_4')

wire n418;
// (7, 8, 'sp4_r_v_b_37')
// (7, 9, 'local_g0_0')
// (7, 9, 'lutff_4/in_2')
// (7, 9, 'sp4_r_v_b_24')
// (7, 10, 'local_g2_0')
// (7, 10, 'local_g3_0')
// (7, 10, 'lutff_6/in_0')
// (7, 10, 'lutff_7/in_0')
// (7, 10, 'neigh_op_tnr_0')
// (7, 10, 'sp4_r_v_b_13')
// (7, 11, 'neigh_op_rgt_0')
// (7, 11, 'sp4_r_v_b_0')
// (7, 12, 'neigh_op_bnr_0')
// (8, 7, 'sp4_v_t_37')
// (8, 8, 'sp4_v_b_37')
// (8, 9, 'local_g2_0')
// (8, 9, 'local_g3_0')
// (8, 9, 'lutff_3/in_0')
// (8, 9, 'lutff_4/in_2')
// (8, 9, 'sp4_v_b_24')
// (8, 10, 'neigh_op_top_0')
// (8, 10, 'sp4_v_b_13')
// (8, 11, 'lutff_0/out')
// (8, 11, 'sp4_v_b_0')
// (8, 12, 'neigh_op_bot_0')
// (9, 10, 'neigh_op_tnl_0')
// (9, 11, 'neigh_op_lft_0')
// (9, 12, 'neigh_op_bnl_0')

wire n419;
// (7, 9, 'local_g2_6')
// (7, 9, 'lutff_1/in_3')
// (7, 9, 'neigh_op_tnr_6')
// (7, 10, 'neigh_op_rgt_6')
// (7, 11, 'neigh_op_bnr_6')
// (8, 9, 'local_g0_6')
// (8, 9, 'local_g1_6')
// (8, 9, 'lutff_3/in_3')
// (8, 9, 'lutff_7/in_2')
// (8, 9, 'neigh_op_top_6')
// (8, 10, 'lutff_6/out')
// (8, 11, 'neigh_op_bot_6')
// (9, 9, 'neigh_op_tnl_6')
// (9, 10, 'neigh_op_lft_6')
// (9, 11, 'neigh_op_bnl_6')

wire n420;
// (7, 9, 'neigh_op_tnr_0')
// (7, 10, 'neigh_op_rgt_0')
// (7, 11, 'neigh_op_bnr_0')
// (8, 9, 'local_g0_0')
// (8, 9, 'local_g1_0')
// (8, 9, 'lutff_5/in_2')
// (8, 9, 'lutff_6/in_2')
// (8, 9, 'neigh_op_top_0')
// (8, 10, 'lutff_0/out')
// (8, 11, 'neigh_op_bot_0')
// (9, 9, 'neigh_op_tnl_0')
// (9, 10, 'neigh_op_lft_0')
// (9, 11, 'neigh_op_bnl_0')

wire n421;
// (7, 9, 'neigh_op_tnr_1')
// (7, 9, 'sp4_r_v_b_47')
// (7, 10, 'neigh_op_rgt_1')
// (7, 10, 'sp4_r_v_b_34')
// (7, 11, 'neigh_op_bnr_1')
// (7, 11, 'sp4_r_v_b_23')
// (7, 12, 'sp4_r_v_b_10')
// (8, 8, 'sp4_v_t_47')
// (8, 9, 'neigh_op_top_1')
// (8, 9, 'sp4_v_b_47')
// (8, 10, 'lutff_1/out')
// (8, 10, 'sp4_h_r_2')
// (8, 10, 'sp4_v_b_34')
// (8, 11, 'local_g0_7')
// (8, 11, 'lutff_0/in_3')
// (8, 11, 'lutff_4/in_3')
// (8, 11, 'neigh_op_bot_1')
// (8, 11, 'sp4_v_b_23')
// (8, 12, 'sp4_v_b_10')
// (9, 9, 'neigh_op_tnl_1')
// (9, 10, 'local_g1_7')
// (9, 10, 'lutff_2/in_0')
// (9, 10, 'neigh_op_lft_1')
// (9, 10, 'sp4_h_r_15')
// (9, 11, 'local_g3_1')
// (9, 11, 'lutff_0/in_0')
// (9, 11, 'lutff_3/in_3')
// (9, 11, 'neigh_op_bnl_1')
// (10, 10, 'sp4_h_r_26')
// (11, 10, 'sp4_h_r_39')
// (12, 10, 'sp4_h_l_39')

wire n422;
// (7, 9, 'neigh_op_tnr_2')
// (7, 10, 'neigh_op_rgt_2')
// (7, 11, 'neigh_op_bnr_2')
// (8, 9, 'neigh_op_top_2')
// (8, 10, 'local_g0_2')
// (8, 10, 'local_g1_2')
// (8, 10, 'lutff_2/out')
// (8, 10, 'lutff_5/in_3')
// (8, 10, 'lutff_7/in_0')
// (8, 11, 'neigh_op_bot_2')
// (9, 9, 'neigh_op_tnl_2')
// (9, 10, 'neigh_op_lft_2')
// (9, 11, 'neigh_op_bnl_2')

wire n423;
// (7, 9, 'neigh_op_tnr_3')
// (7, 10, 'local_g2_3')
// (7, 10, 'lutff_4/in_3')
// (7, 10, 'lutff_5/in_0')
// (7, 10, 'neigh_op_rgt_3')
// (7, 11, 'neigh_op_bnr_3')
// (8, 9, 'neigh_op_top_3')
// (8, 10, 'lutff_3/out')
// (8, 11, 'neigh_op_bot_3')
// (9, 9, 'neigh_op_tnl_3')
// (9, 10, 'local_g1_3')
// (9, 10, 'lutff_6/in_2')
// (9, 10, 'neigh_op_lft_3')
// (9, 11, 'neigh_op_bnl_3')

wire n424;
// (7, 9, 'neigh_op_tnr_4')
// (7, 10, 'local_g2_4')
// (7, 10, 'local_g3_4')
// (7, 10, 'lutff_1/in_3')
// (7, 10, 'lutff_7/in_2')
// (7, 10, 'neigh_op_rgt_4')
// (7, 11, 'neigh_op_bnr_4')
// (8, 9, 'neigh_op_top_4')
// (8, 10, 'lutff_4/out')
// (8, 11, 'neigh_op_bot_4')
// (9, 9, 'neigh_op_tnl_4')
// (9, 10, 'neigh_op_lft_4')
// (9, 11, 'neigh_op_bnl_4')

wire n425;
// (7, 9, 'neigh_op_tnr_5')
// (7, 10, 'neigh_op_rgt_5')
// (7, 11, 'neigh_op_bnr_5')
// (8, 9, 'local_g0_5')
// (8, 9, 'local_g1_5')
// (8, 9, 'lutff_3/in_1')
// (8, 9, 'lutff_4/in_3')
// (8, 9, 'neigh_op_top_5')
// (8, 10, 'lutff_5/out')
// (8, 11, 'neigh_op_bot_5')
// (9, 9, 'neigh_op_tnl_5')
// (9, 10, 'neigh_op_lft_5')
// (9, 11, 'neigh_op_bnl_5')

wire n426;
// (7, 9, 'neigh_op_tnr_7')
// (7, 10, 'neigh_op_rgt_7')
// (7, 11, 'neigh_op_bnr_7')
// (8, 9, 'neigh_op_top_7')
// (8, 10, 'lutff_7/out')
// (8, 11, 'neigh_op_bot_7')
// (9, 9, 'neigh_op_tnl_7')
// (9, 10, 'neigh_op_lft_7')
// (9, 11, 'local_g3_7')
// (9, 11, 'lutff_7/in_3')
// (9, 11, 'neigh_op_bnl_7')

wire n427;
// (7, 10, 'local_g2_2')
// (7, 10, 'local_g3_2')
// (7, 10, 'lutff_1/in_2')
// (7, 10, 'lutff_6/in_1')
// (7, 10, 'lutff_7/in_1')
// (7, 10, 'neigh_op_tnr_2')
// (7, 11, 'neigh_op_rgt_2')
// (7, 12, 'neigh_op_bnr_2')
// (8, 10, 'neigh_op_top_2')
// (8, 11, 'lutff_2/out')
// (8, 12, 'neigh_op_bot_2')
// (9, 10, 'neigh_op_tnl_2')
// (9, 11, 'neigh_op_lft_2')
// (9, 12, 'neigh_op_bnl_2')

wire n428;
// (7, 10, 'neigh_op_tnr_1')
// (7, 11, 'neigh_op_rgt_1')
// (7, 12, 'neigh_op_bnr_1')
// (8, 8, 'sp4_r_v_b_38')
// (8, 9, 'local_g0_3')
// (8, 9, 'local_g1_3')
// (8, 9, 'lutff_5/in_1')
// (8, 9, 'lutff_6/in_1')
// (8, 9, 'lutff_7/in_3')
// (8, 9, 'sp4_r_v_b_27')
// (8, 10, 'neigh_op_top_1')
// (8, 10, 'sp4_r_v_b_14')
// (8, 11, 'lutff_1/out')
// (8, 11, 'sp4_r_v_b_3')
// (8, 12, 'neigh_op_bot_1')
// (9, 7, 'sp4_v_t_38')
// (9, 8, 'sp4_v_b_38')
// (9, 9, 'sp4_v_b_27')
// (9, 10, 'neigh_op_tnl_1')
// (9, 10, 'sp4_v_b_14')
// (9, 11, 'neigh_op_lft_1')
// (9, 11, 'sp4_v_b_3')
// (9, 12, 'neigh_op_bnl_1')

wire n429;
// (7, 10, 'neigh_op_tnr_3')
// (7, 11, 'neigh_op_rgt_3')
// (7, 12, 'neigh_op_bnr_3')
// (8, 10, 'neigh_op_top_3')
// (8, 11, 'local_g0_3')
// (8, 11, 'local_g1_3')
// (8, 11, 'lutff_1/in_2')
// (8, 11, 'lutff_2/in_2')
// (8, 11, 'lutff_3/out')
// (8, 12, 'neigh_op_bot_3')
// (9, 10, 'neigh_op_tnl_3')
// (9, 11, 'neigh_op_lft_3')
// (9, 12, 'neigh_op_bnl_3')

wire n430;
// (7, 10, 'neigh_op_tnr_4')
// (7, 11, 'neigh_op_rgt_4')
// (7, 12, 'neigh_op_bnr_4')
// (8, 8, 'sp4_r_v_b_44')
// (8, 9, 'local_g2_1')
// (8, 9, 'lutff_6/in_3')
// (8, 9, 'sp4_r_v_b_33')
// (8, 10, 'neigh_op_top_4')
// (8, 10, 'sp4_r_v_b_20')
// (8, 11, 'lutff_4/out')
// (8, 11, 'sp4_r_v_b_9')
// (8, 12, 'neigh_op_bot_4')
// (9, 7, 'sp4_v_t_44')
// (9, 8, 'sp4_v_b_44')
// (9, 9, 'sp4_v_b_33')
// (9, 10, 'neigh_op_tnl_4')
// (9, 10, 'sp4_v_b_20')
// (9, 11, 'neigh_op_lft_4')
// (9, 11, 'sp4_v_b_9')
// (9, 12, 'neigh_op_bnl_4')

wire n431;
// (7, 10, 'neigh_op_tnr_6')
// (7, 11, 'neigh_op_rgt_6')
// (7, 12, 'neigh_op_bnr_6')
// (8, 10, 'local_g0_6')
// (8, 10, 'lutff_0/in_0')
// (8, 10, 'lutff_6/in_0')
// (8, 10, 'neigh_op_top_6')
// (8, 11, 'lutff_6/out')
// (8, 12, 'neigh_op_bot_6')
// (9, 10, 'neigh_op_tnl_6')
// (9, 11, 'neigh_op_lft_6')
// (9, 12, 'neigh_op_bnl_6')

wire n432;
// (7, 10, 'neigh_op_tnr_7')
// (7, 11, 'neigh_op_rgt_7')
// (7, 12, 'neigh_op_bnr_7')
// (8, 10, 'local_g0_7')
// (8, 10, 'local_g1_7')
// (8, 10, 'lutff_0/in_2')
// (8, 10, 'lutff_4/in_3')
// (8, 10, 'lutff_5/in_2')
// (8, 10, 'lutff_6/in_3')
// (8, 10, 'neigh_op_top_7')
// (8, 11, 'lutff_7/out')
// (8, 12, 'neigh_op_bot_7')
// (9, 10, 'neigh_op_tnl_7')
// (9, 11, 'neigh_op_lft_7')
// (9, 12, 'neigh_op_bnl_7')

reg n433 = 0;
// (7, 10, 'sp4_r_v_b_40')
// (7, 10, 'sp4_r_v_b_47')
// (7, 11, 'sp4_r_v_b_29')
// (7, 11, 'sp4_r_v_b_34')
// (7, 12, 'local_g0_3')
// (7, 12, 'lutff_5/in_2')
// (7, 12, 'lutff_7/in_0')
// (7, 12, 'sp4_h_r_11')
// (7, 12, 'sp4_r_v_b_16')
// (7, 12, 'sp4_r_v_b_23')
// (7, 13, 'sp4_r_v_b_10')
// (7, 13, 'sp4_r_v_b_5')
// (8, 9, 'sp4_v_t_40')
// (8, 9, 'sp4_v_t_47')
// (8, 10, 'sp4_v_b_40')
// (8, 10, 'sp4_v_b_47')
// (8, 11, 'sp4_v_b_29')
// (8, 11, 'sp4_v_b_34')
// (8, 12, 'local_g0_0')
// (8, 12, 'local_g0_7')
// (8, 12, 'lutff_1/in_2')
// (8, 12, 'lutff_2/in_1')
// (8, 12, 'lutff_5/in_0')
// (8, 12, 'lutff_6/in_0')
// (8, 12, 'sp4_h_r_22')
// (8, 12, 'sp4_v_b_16')
// (8, 12, 'sp4_v_b_23')
// (8, 13, 'local_g0_2')
// (8, 13, 'lutff_7/in_1')
// (8, 13, 'sp4_h_r_5')
// (8, 13, 'sp4_v_b_10')
// (8, 13, 'sp4_v_b_5')
// (9, 12, 'local_g2_3')
// (9, 12, 'lutff_1/in_0')
// (9, 12, 'sp4_h_r_35')
// (9, 13, 'local_g0_0')
// (9, 13, 'lutff_0/in_2')
// (9, 13, 'sp4_h_r_16')
// (10, 12, 'neigh_op_tnr_4')
// (10, 12, 'sp4_h_r_46')
// (10, 13, 'neigh_op_rgt_4')
// (10, 13, 'sp4_h_r_29')
// (10, 13, 'sp4_r_v_b_40')
// (10, 14, 'neigh_op_bnr_4')
// (10, 14, 'sp4_r_v_b_29')
// (10, 15, 'sp4_r_v_b_16')
// (10, 16, 'sp4_r_v_b_5')
// (11, 12, 'local_g1_4')
// (11, 12, 'lutff_1/in_2')
// (11, 12, 'neigh_op_top_4')
// (11, 12, 'sp4_h_l_46')
// (11, 12, 'sp4_v_t_40')
// (11, 13, 'local_g0_4')
// (11, 13, 'lutff_4/in_2')
// (11, 13, 'lutff_4/out')
// (11, 13, 'sp4_h_r_40')
// (11, 13, 'sp4_v_b_40')
// (11, 14, 'neigh_op_bot_4')
// (11, 14, 'sp4_v_b_29')
// (11, 15, 'sp4_v_b_16')
// (11, 16, 'sp4_v_b_5')
// (12, 12, 'neigh_op_tnl_4')
// (12, 13, 'neigh_op_lft_4')
// (12, 13, 'sp4_h_l_40')
// (12, 14, 'neigh_op_bnl_4')

wire n434;
// (7, 11, 'neigh_op_tnr_1')
// (7, 12, 'local_g3_1')
// (7, 12, 'lutff_4/in_2')
// (7, 12, 'neigh_op_rgt_1')
// (7, 13, 'neigh_op_bnr_1')
// (8, 11, 'neigh_op_top_1')
// (8, 12, 'lutff_1/out')
// (8, 13, 'neigh_op_bot_1')
// (9, 11, 'neigh_op_tnl_1')
// (9, 12, 'neigh_op_lft_1')
// (9, 13, 'neigh_op_bnl_1')

wire n435;
// (7, 11, 'neigh_op_tnr_2')
// (7, 12, 'neigh_op_rgt_2')
// (7, 13, 'neigh_op_bnr_2')
// (8, 11, 'neigh_op_top_2')
// (8, 12, 'local_g1_2')
// (8, 12, 'lutff_2/out')
// (8, 12, 'lutff_3/in_0')
// (8, 13, 'neigh_op_bot_2')
// (9, 11, 'neigh_op_tnl_2')
// (9, 12, 'neigh_op_lft_2')
// (9, 13, 'neigh_op_bnl_2')

wire n436;
// (7, 11, 'neigh_op_tnr_3')
// (7, 12, 'local_g2_3')
// (7, 12, 'lutff_3/in_2')
// (7, 12, 'neigh_op_rgt_3')
// (7, 13, 'neigh_op_bnr_3')
// (8, 11, 'neigh_op_top_3')
// (8, 12, 'lutff_3/out')
// (8, 13, 'neigh_op_bot_3')
// (9, 11, 'neigh_op_tnl_3')
// (9, 12, 'neigh_op_lft_3')
// (9, 13, 'neigh_op_bnl_3')

wire n437;
// (7, 11, 'neigh_op_tnr_4')
// (7, 12, 'local_g3_4')
// (7, 12, 'lutff_5/in_0')
// (7, 12, 'lutff_7/in_2')
// (7, 12, 'neigh_op_rgt_4')
// (7, 13, 'neigh_op_bnr_4')
// (8, 11, 'neigh_op_top_4')
// (8, 12, 'lutff_4/out')
// (8, 13, 'neigh_op_bot_4')
// (9, 11, 'neigh_op_tnl_4')
// (9, 12, 'neigh_op_lft_4')
// (9, 13, 'neigh_op_bnl_4')

wire n438;
// (7, 11, 'neigh_op_tnr_5')
// (7, 12, 'neigh_op_rgt_5')
// (7, 13, 'neigh_op_bnr_5')
// (8, 11, 'neigh_op_top_5')
// (8, 12, 'local_g0_5')
// (8, 12, 'lutff_5/out')
// (8, 12, 'lutff_7/in_0')
// (8, 13, 'neigh_op_bot_5')
// (9, 11, 'neigh_op_tnl_5')
// (9, 12, 'neigh_op_lft_5')
// (9, 13, 'neigh_op_bnl_5')

wire n439;
// (7, 11, 'neigh_op_tnr_6')
// (7, 12, 'local_g2_6')
// (7, 12, 'lutff_0/in_2')
// (7, 12, 'neigh_op_rgt_6')
// (7, 13, 'neigh_op_bnr_6')
// (8, 11, 'neigh_op_top_6')
// (8, 12, 'lutff_6/out')
// (8, 13, 'neigh_op_bot_6')
// (9, 11, 'neigh_op_tnl_6')
// (9, 12, 'neigh_op_lft_6')
// (9, 13, 'neigh_op_bnl_6')

wire n440;
// (7, 11, 'neigh_op_tnr_7')
// (7, 12, 'neigh_op_rgt_7')
// (7, 13, 'neigh_op_bnr_7')
// (8, 11, 'neigh_op_top_7')
// (8, 12, 'local_g1_7')
// (8, 12, 'lutff_0/in_2')
// (8, 12, 'lutff_7/out')
// (8, 13, 'neigh_op_bot_7')
// (9, 11, 'neigh_op_tnl_7')
// (9, 12, 'neigh_op_lft_7')
// (9, 13, 'neigh_op_bnl_7')

wire n441;
// (7, 11, 'sp4_r_v_b_38')
// (7, 12, 'local_g1_3')
// (7, 12, 'lutff_1/in_1')
// (7, 12, 'sp4_r_v_b_27')
// (7, 13, 'local_g2_5')
// (7, 13, 'lutff_7/in_0')
// (7, 13, 'neigh_op_tnr_5')
// (7, 13, 'sp4_r_v_b_14')
// (7, 14, 'neigh_op_rgt_5')
// (7, 14, 'sp4_r_v_b_3')
// (7, 15, 'neigh_op_bnr_5')
// (8, 10, 'sp4_v_t_38')
// (8, 11, 'sp4_v_b_38')
// (8, 12, 'sp4_v_b_27')
// (8, 13, 'local_g1_5')
// (8, 13, 'lutff_0/in_0')
// (8, 13, 'lutff_1/in_1')
// (8, 13, 'neigh_op_top_5')
// (8, 13, 'sp4_v_b_14')
// (8, 14, 'lutff_5/out')
// (8, 14, 'sp4_h_r_10')
// (8, 14, 'sp4_v_b_3')
// (8, 15, 'neigh_op_bot_5')
// (9, 13, 'neigh_op_tnl_5')
// (9, 14, 'neigh_op_lft_5')
// (9, 14, 'sp4_h_r_23')
// (9, 15, 'neigh_op_bnl_5')
// (10, 14, 'sp4_h_r_34')
// (11, 14, 'sp4_h_r_47')
// (12, 14, 'sp4_h_l_47')

wire n442;
// (7, 12, 'neigh_op_tnr_0')
// (7, 13, 'neigh_op_rgt_0')
// (7, 14, 'neigh_op_bnr_0')
// (8, 12, 'neigh_op_top_0')
// (8, 13, 'local_g0_0')
// (8, 13, 'lutff_0/out')
// (8, 13, 'lutff_2/in_2')
// (8, 14, 'neigh_op_bot_0')
// (9, 12, 'neigh_op_tnl_0')
// (9, 13, 'neigh_op_lft_0')
// (9, 14, 'neigh_op_bnl_0')

wire n443;
// (7, 12, 'neigh_op_tnr_1')
// (7, 13, 'neigh_op_rgt_1')
// (7, 14, 'neigh_op_bnr_1')
// (8, 12, 'local_g0_1')
// (8, 12, 'lutff_0/in_1')
// (8, 12, 'neigh_op_top_1')
// (8, 13, 'lutff_1/out')
// (8, 14, 'neigh_op_bot_1')
// (9, 12, 'neigh_op_tnl_1')
// (9, 13, 'neigh_op_lft_1')
// (9, 14, 'neigh_op_bnl_1')

wire n444;
// (7, 12, 'neigh_op_tnr_2')
// (7, 13, 'neigh_op_rgt_2')
// (7, 14, 'neigh_op_bnr_2')
// (8, 2, 'sp4_r_v_b_41')
// (8, 3, 'sp4_r_v_b_28')
// (8, 4, 'sp4_r_v_b_17')
// (8, 5, 'sp4_r_v_b_4')
// (8, 6, 'sp4_r_v_b_36')
// (8, 7, 'sp4_r_v_b_25')
// (8, 8, 'sp4_r_v_b_12')
// (8, 9, 'sp4_r_v_b_1')
// (8, 10, 'sp4_r_v_b_40')
// (8, 11, 'sp4_r_v_b_29')
// (8, 12, 'neigh_op_top_2')
// (8, 12, 'sp4_r_v_b_16')
// (8, 13, 'lutff_2/out')
// (8, 13, 'sp4_r_v_b_5')
// (8, 14, 'neigh_op_bot_2')
// (9, 1, 'sp4_v_t_41')
// (9, 2, 'sp4_v_b_41')
// (9, 3, 'sp4_v_b_28')
// (9, 4, 'local_g0_1')
// (9, 4, 'lutff_0/in_1')
// (9, 4, 'sp4_v_b_17')
// (9, 5, 'sp4_h_r_6')
// (9, 5, 'sp4_v_b_4')
// (9, 5, 'sp4_v_t_36')
// (9, 6, 'sp4_v_b_36')
// (9, 7, 'sp4_v_b_25')
// (9, 8, 'sp4_v_b_12')
// (9, 9, 'sp4_v_b_1')
// (9, 9, 'sp4_v_t_40')
// (9, 10, 'sp4_v_b_40')
// (9, 11, 'sp4_v_b_29')
// (9, 12, 'neigh_op_tnl_2')
// (9, 12, 'sp4_v_b_16')
// (9, 13, 'neigh_op_lft_2')
// (9, 13, 'sp4_v_b_5')
// (9, 14, 'neigh_op_bnl_2')
// (10, 2, 'sp4_r_v_b_43')
// (10, 3, 'sp4_r_v_b_30')
// (10, 4, 'sp4_r_v_b_19')
// (10, 5, 'sp4_h_r_19')
// (10, 5, 'sp4_r_v_b_6')
// (11, 1, 'sp4_v_t_43')
// (11, 2, 'sp4_v_b_43')
// (11, 3, 'local_g2_6')
// (11, 3, 'lutff_1/in_1')
// (11, 3, 'sp4_v_b_30')
// (11, 4, 'local_g0_3')
// (11, 4, 'lutff_3/in_2')
// (11, 4, 'sp4_v_b_19')
// (11, 5, 'sp4_h_r_30')
// (11, 5, 'sp4_h_r_6')
// (11, 5, 'sp4_v_b_6')
// (12, 5, 'sp4_h_r_19')
// (12, 5, 'sp4_h_r_43')
// (13, 5, 'span4_horz_19')
// (13, 5, 'span4_horz_43')

wire n445;
// (7, 12, 'neigh_op_tnr_3')
// (7, 13, 'neigh_op_rgt_3')
// (7, 14, 'neigh_op_bnr_3')
// (8, 12, 'neigh_op_top_3')
// (8, 13, 'local_g0_3')
// (8, 13, 'lutff_3/out')
// (8, 13, 'lutff_7/in_2')
// (8, 14, 'neigh_op_bot_3')
// (9, 12, 'neigh_op_tnl_3')
// (9, 13, 'neigh_op_lft_3')
// (9, 14, 'neigh_op_bnl_3')

wire n446;
// (7, 12, 'neigh_op_tnr_5')
// (7, 13, 'neigh_op_rgt_5')
// (7, 14, 'neigh_op_bnr_5')
// (8, 12, 'neigh_op_top_5')
// (8, 13, 'local_g0_5')
// (8, 13, 'lutff_0/in_1')
// (8, 13, 'lutff_1/in_2')
// (8, 13, 'lutff_5/out')
// (8, 14, 'neigh_op_bot_5')
// (9, 12, 'neigh_op_tnl_5')
// (9, 13, 'neigh_op_lft_5')
// (9, 14, 'neigh_op_bnl_5')

wire n447;
// (7, 12, 'neigh_op_tnr_6')
// (7, 13, 'neigh_op_rgt_6')
// (7, 14, 'neigh_op_bnr_6')
// (8, 12, 'neigh_op_top_6')
// (8, 13, 'local_g1_6')
// (8, 13, 'lutff_4/in_1')
// (8, 13, 'lutff_6/out')
// (8, 14, 'neigh_op_bot_6')
// (9, 12, 'neigh_op_tnl_6')
// (9, 13, 'neigh_op_lft_6')
// (9, 14, 'neigh_op_bnl_6')

wire n448;
// (7, 12, 'neigh_op_tnr_7')
// (7, 13, 'neigh_op_rgt_7')
// (7, 14, 'neigh_op_bnr_7')
// (8, 12, 'neigh_op_top_7')
// (8, 13, 'local_g0_7')
// (8, 13, 'lutff_2/in_1')
// (8, 13, 'lutff_7/out')
// (8, 14, 'neigh_op_bot_7')
// (9, 12, 'neigh_op_tnl_7')
// (9, 13, 'neigh_op_lft_7')
// (9, 14, 'neigh_op_bnl_7')

wire n449;
// (7, 13, 'local_g2_0')
// (7, 13, 'lutff_4/in_0')
// (7, 13, 'neigh_op_tnr_0')
// (7, 14, 'neigh_op_rgt_0')
// (7, 15, 'neigh_op_bnr_0')
// (8, 11, 'sp4_r_v_b_36')
// (8, 12, 'sp4_r_v_b_25')
// (8, 13, 'local_g2_4')
// (8, 13, 'lutff_5/in_3')
// (8, 13, 'neigh_op_top_0')
// (8, 13, 'sp4_r_v_b_12')
// (8, 14, 'lutff_0/out')
// (8, 14, 'sp4_r_v_b_1')
// (8, 15, 'neigh_op_bot_0')
// (9, 10, 'sp4_v_t_36')
// (9, 11, 'sp4_v_b_36')
// (9, 12, 'sp4_v_b_25')
// (9, 13, 'neigh_op_tnl_0')
// (9, 13, 'sp4_v_b_12')
// (9, 14, 'neigh_op_lft_0')
// (9, 14, 'sp4_v_b_1')
// (9, 15, 'neigh_op_bnl_0')

wire n450;
// (7, 13, 'local_g3_4')
// (7, 13, 'lutff_6/in_1')
// (7, 13, 'neigh_op_tnr_4')
// (7, 14, 'neigh_op_rgt_4')
// (7, 15, 'neigh_op_bnr_4')
// (8, 13, 'local_g1_4')
// (8, 13, 'lutff_0/in_3')
// (8, 13, 'lutff_6/in_1')
// (8, 13, 'neigh_op_top_4')
// (8, 14, 'lutff_4/out')
// (8, 15, 'neigh_op_bot_4')
// (9, 13, 'neigh_op_tnl_4')
// (9, 14, 'neigh_op_lft_4')
// (9, 15, 'neigh_op_bnl_4')

wire n451;
// (7, 13, 'neigh_op_tnr_1')
// (7, 14, 'neigh_op_rgt_1')
// (7, 15, 'neigh_op_bnr_1')
// (8, 13, 'neigh_op_top_1')
// (8, 14, 'local_g0_1')
// (8, 14, 'local_g1_1')
// (8, 14, 'lutff_1/out')
// (8, 14, 'lutff_4/in_0')
// (8, 14, 'lutff_5/in_0')
// (8, 14, 'lutff_6/in_0')
// (8, 14, 'lutff_7/in_0')
// (8, 15, 'neigh_op_bot_1')
// (9, 13, 'neigh_op_tnl_1')
// (9, 14, 'neigh_op_lft_1')
// (9, 15, 'neigh_op_bnl_1')

wire n452;
// (7, 13, 'neigh_op_tnr_2')
// (7, 14, 'neigh_op_rgt_2')
// (7, 15, 'neigh_op_bnr_2')
// (8, 13, 'neigh_op_top_2')
// (8, 14, 'local_g0_2')
// (8, 14, 'local_g1_2')
// (8, 14, 'lutff_2/out')
// (8, 14, 'lutff_4/in_1')
// (8, 14, 'lutff_5/in_2')
// (8, 14, 'lutff_6/in_1')
// (8, 14, 'lutff_7/in_1')
// (8, 15, 'neigh_op_bot_2')
// (9, 13, 'neigh_op_tnl_2')
// (9, 14, 'neigh_op_lft_2')
// (9, 15, 'neigh_op_bnl_2')

wire n453;
// (7, 13, 'neigh_op_tnr_3')
// (7, 14, 'neigh_op_rgt_3')
// (7, 15, 'local_g0_3')
// (7, 15, 'local_g1_3')
// (7, 15, 'lutff_0/in_2')
// (7, 15, 'lutff_4/in_2')
// (7, 15, 'lutff_6/in_1')
// (7, 15, 'neigh_op_bnr_3')
// (8, 13, 'neigh_op_top_3')
// (8, 14, 'lutff_3/out')
// (8, 15, 'neigh_op_bot_3')
// (9, 13, 'neigh_op_tnl_3')
// (9, 14, 'neigh_op_lft_3')
// (9, 15, 'neigh_op_bnl_3')

wire n454;
// (7, 13, 'neigh_op_tnr_6')
// (7, 14, 'neigh_op_rgt_6')
// (7, 15, 'neigh_op_bnr_6')
// (8, 12, 'sp4_r_v_b_37')
// (8, 13, 'local_g1_0')
// (8, 13, 'lutff_6/in_3')
// (8, 13, 'neigh_op_top_6')
// (8, 13, 'sp4_r_v_b_24')
// (8, 14, 'lutff_6/out')
// (8, 14, 'sp4_r_v_b_13')
// (8, 15, 'neigh_op_bot_6')
// (8, 15, 'sp4_r_v_b_0')
// (9, 11, 'sp4_v_t_37')
// (9, 12, 'sp4_v_b_37')
// (9, 13, 'neigh_op_tnl_6')
// (9, 13, 'sp4_v_b_24')
// (9, 14, 'neigh_op_lft_6')
// (9, 14, 'sp4_v_b_13')
// (9, 15, 'neigh_op_bnl_6')
// (9, 15, 'sp4_v_b_0')

reg n455 = 0;
// (7, 13, 'sp4_r_v_b_45')
// (7, 14, 'sp4_r_v_b_32')
// (7, 15, 'sp4_r_v_b_21')
// (7, 16, 'sp4_r_v_b_8')
// (8, 12, 'local_g1_0')
// (8, 12, 'local_g1_1')
// (8, 12, 'lutff_1/in_0')
// (8, 12, 'lutff_2/in_0')
// (8, 12, 'lutff_4/in_3')
// (8, 12, 'lutff_5/in_3')
// (8, 12, 'lutff_6/in_3')
// (8, 12, 'sp4_h_r_1')
// (8, 12, 'sp4_h_r_8')
// (8, 12, 'sp4_v_t_45')
// (8, 13, 'local_g0_1')
// (8, 13, 'lutff_3/in_2')
// (8, 13, 'sp4_h_r_9')
// (8, 13, 'sp4_v_b_45')
// (8, 14, 'sp4_v_b_32')
// (8, 15, 'sp4_v_b_21')
// (8, 16, 'sp4_v_b_8')
// (9, 12, 'local_g1_5')
// (9, 12, 'lutff_1/in_1')
// (9, 12, 'sp4_h_r_12')
// (9, 12, 'sp4_h_r_21')
// (9, 13, 'local_g0_4')
// (9, 13, 'lutff_2/in_2')
// (9, 13, 'sp4_h_r_20')
// (10, 12, 'neigh_op_tnr_6')
// (10, 12, 'sp4_h_r_25')
// (10, 12, 'sp4_h_r_32')
// (10, 13, 'neigh_op_rgt_6')
// (10, 13, 'sp4_h_r_33')
// (10, 14, 'neigh_op_bnr_6')
// (11, 12, 'local_g0_6')
// (11, 12, 'lutff_1/in_1')
// (11, 12, 'neigh_op_top_6')
// (11, 12, 'sp4_h_r_36')
// (11, 12, 'sp4_h_r_45')
// (11, 13, 'local_g0_6')
// (11, 13, 'lutff_6/in_2')
// (11, 13, 'lutff_6/out')
// (11, 13, 'sp4_h_r_44')
// (11, 13, 'sp4_r_v_b_45')
// (11, 14, 'neigh_op_bot_6')
// (11, 14, 'sp4_r_v_b_32')
// (11, 15, 'sp4_r_v_b_21')
// (11, 16, 'sp4_r_v_b_8')
// (12, 12, 'neigh_op_tnl_6')
// (12, 12, 'sp4_h_l_36')
// (12, 12, 'sp4_h_l_45')
// (12, 12, 'sp4_v_t_45')
// (12, 13, 'neigh_op_lft_6')
// (12, 13, 'sp4_h_l_44')
// (12, 13, 'sp4_v_b_45')
// (12, 14, 'neigh_op_bnl_6')
// (12, 14, 'sp4_v_b_32')
// (12, 15, 'sp4_v_b_21')
// (12, 16, 'sp4_v_b_8')

reg \d_out[1] = 0 ;
// (8, 1, 'sp4_r_v_b_34')
// (8, 2, 'sp4_r_v_b_23')
// (8, 3, 'sp4_r_v_b_10')
// (9, 0, 'io_0/D_OUT_0')
// (9, 0, 'io_0/PAD')
// (9, 0, 'local_g0_2')
// (9, 0, 'span4_vert_34')
// (9, 1, 'sp4_v_b_34')
// (9, 2, 'sp4_v_b_23')
// (9, 3, 'sp4_h_r_10')
// (9, 3, 'sp4_v_b_10')
// (10, 2, 'neigh_op_tnr_1')
// (10, 3, 'neigh_op_rgt_1')
// (10, 3, 'sp4_h_r_23')
// (10, 4, 'neigh_op_bnr_1')
// (11, 2, 'neigh_op_top_1')
// (11, 3, 'lutff_1/out')
// (11, 3, 'sp4_h_r_34')
// (11, 4, 'neigh_op_bot_1')
// (12, 2, 'neigh_op_tnl_1')
// (12, 3, 'neigh_op_lft_1')
// (12, 3, 'sp4_h_r_47')
// (12, 4, 'neigh_op_bnl_1')
// (13, 3, 'span4_horz_47')

reg n457 = 0;
// (8, 2, 'neigh_op_tnr_3')
// (8, 3, 'neigh_op_rgt_3')
// (8, 4, 'neigh_op_bnr_3')
// (9, 2, 'neigh_op_top_3')
// (9, 3, 'local_g1_3')
// (9, 3, 'lutff_3/out')
// (9, 3, 'lutff_6/in_0')
// (9, 4, 'neigh_op_bot_3')
// (10, 2, 'neigh_op_tnl_3')
// (10, 3, 'neigh_op_lft_3')
// (10, 4, 'neigh_op_bnl_3')

reg n458 = 0;
// (8, 2, 'neigh_op_tnr_4')
// (8, 3, 'neigh_op_rgt_4')
// (8, 4, 'neigh_op_bnr_4')
// (9, 2, 'neigh_op_top_4')
// (9, 3, 'local_g1_4')
// (9, 3, 'lutff_4/out')
// (9, 3, 'lutff_5/in_0')
// (9, 4, 'neigh_op_bot_4')
// (10, 2, 'neigh_op_tnl_4')
// (10, 3, 'neigh_op_lft_4')
// (10, 4, 'neigh_op_bnl_4')

reg n459 = 0;
// (8, 2, 'neigh_op_tnr_5')
// (8, 3, 'neigh_op_rgt_5')
// (8, 4, 'neigh_op_bnr_5')
// (9, 2, 'neigh_op_top_5')
// (9, 3, 'local_g0_5')
// (9, 3, 'lutff_3/in_0')
// (9, 3, 'lutff_5/out')
// (9, 4, 'neigh_op_bot_5')
// (10, 2, 'neigh_op_tnl_5')
// (10, 3, 'neigh_op_lft_5')
// (10, 4, 'neigh_op_bnl_5')

reg n460 = 0;
// (8, 2, 'neigh_op_tnr_6')
// (8, 3, 'local_g2_6')
// (8, 3, 'local_g3_6')
// (8, 3, 'lutff_1/in_1')
// (8, 3, 'lutff_3/in_2')
// (8, 3, 'lutff_6/in_0')
// (8, 3, 'neigh_op_rgt_6')
// (8, 4, 'neigh_op_bnr_6')
// (9, 2, 'neigh_op_top_6')
// (9, 3, 'local_g0_6')
// (9, 3, 'lutff_4/in_0')
// (9, 3, 'lutff_6/out')
// (9, 4, 'neigh_op_bot_6')
// (10, 2, 'neigh_op_tnl_6')
// (10, 3, 'neigh_op_lft_6')
// (10, 4, 'neigh_op_bnl_6')

reg n461 = 0;
// (8, 3, 'neigh_op_tnr_0')
// (8, 4, 'neigh_op_rgt_0')
// (8, 5, 'neigh_op_bnr_0')
// (9, 3, 'neigh_op_top_0')
// (9, 4, 'local_g1_0')
// (9, 4, 'lutff_0/out')
// (9, 4, 'lutff_1/in_0')
// (9, 5, 'neigh_op_bot_0')
// (10, 3, 'neigh_op_tnl_0')
// (10, 4, 'neigh_op_lft_0')
// (10, 5, 'neigh_op_bnl_0')

reg n462 = 0;
// (8, 3, 'neigh_op_tnr_1')
// (8, 4, 'neigh_op_rgt_1')
// (8, 5, 'neigh_op_bnr_1')
// (9, 3, 'neigh_op_top_1')
// (9, 4, 'local_g1_1')
// (9, 4, 'lutff_1/out')
// (9, 4, 'lutff_6/in_0')
// (9, 5, 'neigh_op_bot_1')
// (10, 3, 'neigh_op_tnl_1')
// (10, 4, 'neigh_op_lft_1')
// (10, 5, 'neigh_op_bnl_1')

reg n463 = 0;
// (8, 3, 'neigh_op_tnr_4')
// (8, 4, 'neigh_op_rgt_4')
// (8, 5, 'neigh_op_bnr_4')
// (9, 3, 'neigh_op_top_4')
// (9, 4, 'local_g1_4')
// (9, 4, 'lutff_0/in_3')
// (9, 4, 'lutff_4/out')
// (9, 5, 'neigh_op_bot_4')
// (10, 3, 'neigh_op_tnl_4')
// (10, 4, 'neigh_op_lft_4')
// (10, 5, 'neigh_op_bnl_4')

reg n464 = 0;
// (8, 3, 'neigh_op_tnr_6')
// (8, 4, 'neigh_op_rgt_6')
// (8, 5, 'neigh_op_bnr_6')
// (9, 3, 'neigh_op_top_6')
// (9, 4, 'local_g1_6')
// (9, 4, 'lutff_6/out')
// (9, 4, 'lutff_7/in_0')
// (9, 5, 'neigh_op_bot_6')
// (10, 3, 'neigh_op_tnl_6')
// (10, 4, 'neigh_op_lft_6')
// (10, 5, 'neigh_op_bnl_6')

reg n465 = 0;
// (8, 4, 'neigh_op_tnr_0')
// (8, 5, 'neigh_op_rgt_0')
// (8, 6, 'neigh_op_bnr_0')
// (9, 4, 'local_g0_0')
// (9, 4, 'lutff_4/in_0')
// (9, 4, 'neigh_op_top_0')
// (9, 5, 'lutff_0/out')
// (9, 6, 'neigh_op_bot_0')
// (10, 4, 'neigh_op_tnl_0')
// (10, 5, 'neigh_op_lft_0')
// (10, 6, 'neigh_op_bnl_0')

reg n466 = 0;
// (8, 4, 'neigh_op_tnr_1')
// (8, 5, 'neigh_op_rgt_1')
// (8, 6, 'neigh_op_bnr_1')
// (9, 4, 'neigh_op_top_1')
// (9, 5, 'local_g1_1')
// (9, 5, 'lutff_1/out')
// (9, 5, 'lutff_4/in_0')
// (9, 6, 'neigh_op_bot_1')
// (10, 4, 'neigh_op_tnl_1')
// (10, 5, 'neigh_op_lft_1')
// (10, 6, 'neigh_op_bnl_1')

reg n467 = 0;
// (8, 4, 'neigh_op_tnr_2')
// (8, 5, 'neigh_op_rgt_2')
// (8, 6, 'neigh_op_bnr_2')
// (9, 4, 'neigh_op_top_2')
// (9, 5, 'lutff_2/out')
// (9, 6, 'local_g0_2')
// (9, 6, 'lutff_2/in_0')
// (9, 6, 'neigh_op_bot_2')
// (10, 4, 'neigh_op_tnl_2')
// (10, 5, 'neigh_op_lft_2')
// (10, 6, 'neigh_op_bnl_2')

reg n468 = 0;
// (8, 4, 'neigh_op_tnr_3')
// (8, 5, 'neigh_op_rgt_3')
// (8, 6, 'neigh_op_bnr_3')
// (9, 4, 'neigh_op_top_3')
// (9, 5, 'local_g1_3')
// (9, 5, 'lutff_0/in_0')
// (9, 5, 'lutff_3/out')
// (9, 6, 'neigh_op_bot_3')
// (10, 4, 'neigh_op_tnl_3')
// (10, 5, 'neigh_op_lft_3')
// (10, 6, 'neigh_op_bnl_3')

reg n469 = 0;
// (8, 4, 'neigh_op_tnr_4')
// (8, 5, 'neigh_op_rgt_4')
// (8, 6, 'neigh_op_bnr_4')
// (9, 4, 'neigh_op_top_4')
// (9, 5, 'local_g0_4')
// (9, 5, 'lutff_4/out')
// (9, 5, 'lutff_6/in_0')
// (9, 6, 'neigh_op_bot_4')
// (10, 4, 'neigh_op_tnl_4')
// (10, 5, 'neigh_op_lft_4')
// (10, 6, 'neigh_op_bnl_4')

reg n470 = 0;
// (8, 4, 'neigh_op_tnr_5')
// (8, 5, 'neigh_op_rgt_5')
// (8, 6, 'neigh_op_bnr_5')
// (9, 4, 'neigh_op_top_5')
// (9, 5, 'local_g2_5')
// (9, 5, 'lutff_3/in_0')
// (9, 5, 'lutff_5/out')
// (9, 6, 'neigh_op_bot_5')
// (10, 4, 'neigh_op_tnl_5')
// (10, 5, 'neigh_op_lft_5')
// (10, 6, 'neigh_op_bnl_5')

reg n471 = 0;
// (8, 4, 'neigh_op_tnr_6')
// (8, 5, 'neigh_op_rgt_6')
// (8, 6, 'neigh_op_bnr_6')
// (9, 4, 'neigh_op_top_6')
// (9, 5, 'local_g1_6')
// (9, 5, 'lutff_5/in_0')
// (9, 5, 'lutff_6/out')
// (9, 6, 'neigh_op_bot_6')
// (10, 4, 'neigh_op_tnl_6')
// (10, 5, 'neigh_op_lft_6')
// (10, 6, 'neigh_op_bnl_6')

wire n472;
// (8, 5, 'neigh_op_tnr_0')
// (8, 6, 'neigh_op_rgt_0')
// (8, 7, 'neigh_op_bnr_0')
// (9, 5, 'neigh_op_top_0')
// (9, 6, 'lutff_0/out')
// (9, 7, 'local_g0_0')
// (9, 7, 'lutff_0/in_0')
// (9, 7, 'neigh_op_bot_0')
// (10, 5, 'neigh_op_tnl_0')
// (10, 6, 'neigh_op_lft_0')
// (10, 7, 'neigh_op_bnl_0')

reg n473 = 0;
// (8, 5, 'neigh_op_tnr_2')
// (8, 6, 'neigh_op_rgt_2')
// (8, 7, 'neigh_op_bnr_2')
// (9, 5, 'neigh_op_top_2')
// (9, 6, 'local_g1_2')
// (9, 6, 'lutff_2/out')
// (9, 6, 'lutff_7/in_0')
// (9, 7, 'neigh_op_bot_2')
// (10, 5, 'neigh_op_tnl_2')
// (10, 6, 'neigh_op_lft_2')
// (10, 7, 'neigh_op_bnl_2')

reg n474 = 0;
// (8, 5, 'neigh_op_tnr_4')
// (8, 6, 'neigh_op_rgt_4')
// (8, 7, 'neigh_op_bnr_4')
// (9, 5, 'neigh_op_top_4')
// (9, 6, 'local_g1_4')
// (9, 6, 'lutff_1/in_0')
// (9, 6, 'lutff_4/out')
// (9, 7, 'neigh_op_bot_4')
// (10, 5, 'neigh_op_tnl_4')
// (10, 6, 'neigh_op_lft_4')
// (10, 7, 'neigh_op_bnl_4')

reg n475 = 0;
// (8, 5, 'neigh_op_tnr_5')
// (8, 6, 'neigh_op_rgt_5')
// (8, 7, 'neigh_op_bnr_5')
// (9, 5, 'local_g0_5')
// (9, 5, 'lutff_1/in_0')
// (9, 5, 'neigh_op_top_5')
// (9, 6, 'lutff_5/out')
// (9, 7, 'neigh_op_bot_5')
// (10, 5, 'neigh_op_tnl_5')
// (10, 6, 'neigh_op_lft_5')
// (10, 7, 'neigh_op_bnl_5')

reg n476 = 0;
// (8, 5, 'neigh_op_tnr_6')
// (8, 6, 'neigh_op_rgt_6')
// (8, 7, 'neigh_op_bnr_6')
// (9, 5, 'local_g0_6')
// (9, 5, 'lutff_2/in_0')
// (9, 5, 'neigh_op_top_6')
// (9, 6, 'lutff_6/out')
// (9, 7, 'neigh_op_bot_6')
// (10, 5, 'neigh_op_tnl_6')
// (10, 6, 'neigh_op_lft_6')
// (10, 7, 'neigh_op_bnl_6')

reg n477 = 0;
// (8, 5, 'neigh_op_tnr_7')
// (8, 6, 'neigh_op_rgt_7')
// (8, 7, 'neigh_op_bnr_7')
// (9, 5, 'neigh_op_top_7')
// (9, 6, 'local_g0_7')
// (9, 6, 'local_g1_7')
// (9, 6, 'lutff_0/in_1')
// (9, 6, 'lutff_3/in_0')
// (9, 6, 'lutff_4/in_2')
// (9, 6, 'lutff_6/in_0')
// (9, 6, 'lutff_7/out')
// (9, 7, 'neigh_op_bot_7')
// (10, 5, 'neigh_op_tnl_7')
// (10, 6, 'neigh_op_lft_7')
// (10, 7, 'neigh_op_bnl_7')

wire n478;
// (8, 6, 'neigh_op_tnr_0')
// (8, 6, 'sp4_r_v_b_45')
// (8, 7, 'neigh_op_rgt_0')
// (8, 7, 'sp4_r_v_b_32')
// (8, 8, 'neigh_op_bnr_0')
// (8, 8, 'sp4_r_v_b_21')
// (8, 9, 'sp4_r_v_b_8')
// (8, 10, 'sp4_r_v_b_41')
// (8, 11, 'sp4_r_v_b_28')
// (8, 12, 'sp4_r_v_b_17')
// (8, 13, 'sp4_r_v_b_4')
// (9, 5, 'sp4_v_t_45')
// (9, 6, 'neigh_op_top_0')
// (9, 6, 'sp4_v_b_45')
// (9, 7, 'lutff_0/out')
// (9, 7, 'sp4_v_b_32')
// (9, 8, 'neigh_op_bot_0')
// (9, 8, 'sp4_v_b_21')
// (9, 9, 'local_g0_0')
// (9, 9, 'local_g1_0')
// (9, 9, 'lutff_1/in_2')
// (9, 9, 'lutff_4/in_2')
// (9, 9, 'sp4_v_b_8')
// (9, 9, 'sp4_v_t_41')
// (9, 10, 'local_g2_1')
// (9, 10, 'local_g3_1')
// (9, 10, 'lutff_1/in_2')
// (9, 10, 'lutff_3/in_3')
// (9, 10, 'lutff_4/in_2')
// (9, 10, 'sp4_v_b_41')
// (9, 11, 'sp4_v_b_28')
// (9, 12, 'sp4_v_b_17')
// (9, 13, 'sp4_v_b_4')
// (10, 6, 'neigh_op_tnl_0')
// (10, 7, 'neigh_op_lft_0')
// (10, 8, 'neigh_op_bnl_0')

wire n479;
// (8, 6, 'neigh_op_tnr_1')
// (8, 7, 'neigh_op_rgt_1')
// (8, 8, 'neigh_op_bnr_1')
// (9, 6, 'neigh_op_top_1')
// (9, 7, 'local_g2_1')
// (9, 7, 'lutff_1/out')
// (9, 7, 'lutff_2/in_3')
// (9, 8, 'neigh_op_bot_1')
// (10, 6, 'neigh_op_tnl_1')
// (10, 7, 'neigh_op_lft_1')
// (10, 8, 'neigh_op_bnl_1')

wire n480;
// (8, 6, 'neigh_op_tnr_2')
// (8, 7, 'neigh_op_rgt_2')
// (8, 7, 'sp4_r_v_b_36')
// (8, 8, 'neigh_op_bnr_2')
// (8, 8, 'sp4_r_v_b_25')
// (8, 9, 'sp4_r_v_b_12')
// (8, 10, 'sp4_r_v_b_1')
// (9, 6, 'neigh_op_top_2')
// (9, 6, 'sp4_v_t_36')
// (9, 7, 'lutff_2/out')
// (9, 7, 'sp4_v_b_36')
// (9, 8, 'neigh_op_bot_2')
// (9, 8, 'sp4_v_b_25')
// (9, 9, 'local_g0_4')
// (9, 9, 'local_g1_4')
// (9, 9, 'lutff_0/in_3')
// (9, 9, 'lutff_5/in_3')
// (9, 9, 'sp4_v_b_12')
// (9, 10, 'sp4_v_b_1')
// (10, 6, 'neigh_op_tnl_2')
// (10, 7, 'neigh_op_lft_2')
// (10, 8, 'neigh_op_bnl_2')

reg n481 = 0;
// (8, 6, 'neigh_op_tnr_5')
// (8, 7, 'neigh_op_rgt_5')
// (8, 7, 'sp12_h_r_1')
// (8, 8, 'neigh_op_bnr_5')
// (9, 6, 'neigh_op_top_5')
// (9, 7, 'lutff_5/out')
// (9, 7, 'sp12_h_r_2')
// (9, 8, 'neigh_op_bot_5')
// (10, 6, 'neigh_op_tnl_5')
// (10, 7, 'neigh_op_lft_5')
// (10, 7, 'sp12_h_r_5')
// (10, 8, 'neigh_op_bnl_5')
// (11, 7, 'local_g0_6')
// (11, 7, 'lutff_2/in_0')
// (11, 7, 'sp12_h_r_6')
// (12, 7, 'sp12_h_r_9')
// (13, 7, 'span12_horz_9')

reg n482 = 0;
// (8, 6, 'neigh_op_tnr_6')
// (8, 7, 'neigh_op_rgt_6')
// (8, 8, 'neigh_op_bnr_6')
// (9, 6, 'neigh_op_top_6')
// (9, 6, 'sp4_r_v_b_40')
// (9, 7, 'local_g1_5')
// (9, 7, 'local_g1_6')
// (9, 7, 'lutff_1/in_0')
// (9, 7, 'lutff_5/in_1')
// (9, 7, 'lutff_6/out')
// (9, 7, 'sp4_r_v_b_29')
// (9, 8, 'neigh_op_bot_6')
// (9, 8, 'sp4_r_v_b_16')
// (9, 9, 'sp4_r_v_b_5')
// (10, 5, 'sp4_v_t_40')
// (10, 6, 'neigh_op_tnl_6')
// (10, 6, 'sp4_v_b_40')
// (10, 7, 'neigh_op_lft_6')
// (10, 7, 'sp4_v_b_29')
// (10, 8, 'neigh_op_bnl_6')
// (10, 8, 'sp4_v_b_16')
// (10, 9, 'sp4_v_b_5')

reg n483 = 0;
// (8, 6, 'neigh_op_tnr_7')
// (8, 7, 'neigh_op_rgt_7')
// (8, 8, 'neigh_op_bnr_7')
// (9, 6, 'neigh_op_top_7')
// (9, 7, 'local_g1_7')
// (9, 7, 'lutff_6/in_0')
// (9, 7, 'lutff_7/out')
// (9, 8, 'neigh_op_bot_7')
// (10, 6, 'neigh_op_tnl_7')
// (10, 7, 'neigh_op_lft_7')
// (10, 8, 'neigh_op_bnl_7')

reg n484 = 0;
// (8, 6, 'sp4_h_r_11')
// (9, 6, 'local_g0_6')
// (9, 6, 'lutff_3/in_1')
// (9, 6, 'sp4_h_r_22')
// (10, 5, 'neigh_op_tnr_7')
// (10, 6, 'neigh_op_rgt_7')
// (10, 6, 'sp4_h_r_35')
// (10, 7, 'neigh_op_bnr_7')
// (11, 5, 'neigh_op_top_7')
// (11, 6, 'local_g0_7')
// (11, 6, 'lutff_0/in_1')
// (11, 6, 'lutff_7/out')
// (11, 6, 'sp4_h_r_46')
// (11, 7, 'neigh_op_bot_7')
// (12, 5, 'neigh_op_tnl_7')
// (12, 6, 'neigh_op_lft_7')
// (12, 6, 'sp4_h_l_46')
// (12, 7, 'neigh_op_bnl_7')

reg n485 = 0;
// (8, 6, 'sp4_h_r_5')
// (9, 6, 'local_g1_0')
// (9, 6, 'lutff_6/in_1')
// (9, 6, 'sp4_h_r_16')
// (10, 5, 'neigh_op_tnr_4')
// (10, 6, 'neigh_op_rgt_4')
// (10, 6, 'sp4_h_r_29')
// (10, 7, 'neigh_op_bnr_4')
// (11, 5, 'neigh_op_top_4')
// (11, 6, 'local_g0_4')
// (11, 6, 'lutff_0/in_0')
// (11, 6, 'lutff_4/out')
// (11, 6, 'sp4_h_r_40')
// (11, 7, 'neigh_op_bot_4')
// (12, 5, 'neigh_op_tnl_4')
// (12, 6, 'neigh_op_lft_4')
// (12, 6, 'sp4_h_l_40')
// (12, 7, 'neigh_op_bnl_4')

reg n486 = 0;
// (8, 7, 'local_g0_1')
// (8, 7, 'lutff_0/in_1')
// (8, 7, 'sp4_h_r_1')
// (9, 7, 'sp4_h_r_12')
// (10, 6, 'neigh_op_tnr_0')
// (10, 7, 'neigh_op_rgt_0')
// (10, 7, 'sp4_h_r_25')
// (10, 8, 'neigh_op_bnr_0')
// (11, 4, 'sp4_r_v_b_36')
// (11, 5, 'sp4_r_v_b_25')
// (11, 6, 'neigh_op_top_0')
// (11, 6, 'sp4_r_v_b_12')
// (11, 7, 'lutff_0/out')
// (11, 7, 'sp4_h_r_36')
// (11, 7, 'sp4_r_v_b_1')
// (11, 8, 'neigh_op_bot_0')
// (12, 3, 'sp4_v_t_36')
// (12, 4, 'sp4_v_b_36')
// (12, 5, 'sp4_v_b_25')
// (12, 6, 'neigh_op_tnl_0')
// (12, 6, 'sp4_v_b_12')
// (12, 7, 'neigh_op_lft_0')
// (12, 7, 'sp4_h_l_36')
// (12, 7, 'sp4_v_b_1')
// (12, 8, 'neigh_op_bnl_0')

reg n487 = 0;
// (8, 7, 'neigh_op_tnr_0')
// (8, 8, 'neigh_op_rgt_0')
// (8, 9, 'neigh_op_bnr_0')
// (9, 7, 'neigh_op_top_0')
// (9, 8, 'local_g1_0')
// (9, 8, 'lutff_0/out')
// (9, 8, 'lutff_1/in_0')
// (9, 9, 'neigh_op_bot_0')
// (10, 7, 'neigh_op_tnl_0')
// (10, 8, 'neigh_op_lft_0')
// (10, 9, 'neigh_op_bnl_0')

reg n488 = 0;
// (8, 7, 'neigh_op_tnr_1')
// (8, 8, 'neigh_op_rgt_1')
// (8, 9, 'neigh_op_bnr_1')
// (9, 7, 'neigh_op_top_1')
// (9, 8, 'local_g1_1')
// (9, 8, 'lutff_1/out')
// (9, 8, 'lutff_4/in_0')
// (9, 9, 'neigh_op_bot_1')
// (10, 7, 'neigh_op_tnl_1')
// (10, 8, 'neigh_op_lft_1')
// (10, 9, 'neigh_op_bnl_1')

reg n489 = 0;
// (8, 7, 'neigh_op_tnr_2')
// (8, 8, 'neigh_op_rgt_2')
// (8, 9, 'neigh_op_bnr_2')
// (9, 7, 'neigh_op_top_2')
// (9, 8, 'local_g1_2')
// (9, 8, 'lutff_2/out')
// (9, 8, 'lutff_5/in_0')
// (9, 9, 'neigh_op_bot_2')
// (10, 7, 'neigh_op_tnl_2')
// (10, 8, 'neigh_op_lft_2')
// (10, 9, 'neigh_op_bnl_2')

reg n490 = 0;
// (8, 7, 'neigh_op_tnr_4')
// (8, 8, 'neigh_op_rgt_4')
// (8, 9, 'neigh_op_bnr_4')
// (9, 7, 'neigh_op_top_4')
// (9, 8, 'local_g0_4')
// (9, 8, 'lutff_2/in_0')
// (9, 8, 'lutff_4/out')
// (9, 9, 'neigh_op_bot_4')
// (10, 7, 'neigh_op_tnl_4')
// (10, 8, 'neigh_op_lft_4')
// (10, 9, 'neigh_op_bnl_4')

reg n491 = 0;
// (8, 7, 'neigh_op_tnr_5')
// (8, 8, 'neigh_op_rgt_5')
// (8, 9, 'neigh_op_bnr_5')
// (9, 7, 'neigh_op_top_5')
// (9, 8, 'local_g0_5')
// (9, 8, 'lutff_5/out')
// (9, 8, 'lutff_7/in_0')
// (9, 9, 'neigh_op_bot_5')
// (10, 7, 'neigh_op_tnl_5')
// (10, 8, 'neigh_op_lft_5')
// (10, 9, 'neigh_op_bnl_5')

wire n492;
// (8, 7, 'sp4_h_r_3')
// (9, 7, 'local_g0_6')
// (9, 7, 'lutff_2/in_0')
// (9, 7, 'sp4_h_r_14')
// (10, 7, 'sp4_h_r_27')
// (10, 8, 'neigh_op_tnr_0')
// (10, 9, 'neigh_op_rgt_0')
// (10, 10, 'neigh_op_bnr_0')
// (11, 6, 'sp4_r_v_b_36')
// (11, 7, 'local_g0_1')
// (11, 7, 'lutff_4/in_1')
// (11, 7, 'sp4_h_r_38')
// (11, 7, 'sp4_r_v_b_25')
// (11, 8, 'neigh_op_top_0')
// (11, 8, 'sp4_r_v_b_12')
// (11, 8, 'sp4_r_v_b_44')
// (11, 9, 'lutff_0/out')
// (11, 9, 'sp4_r_v_b_1')
// (11, 9, 'sp4_r_v_b_33')
// (11, 10, 'neigh_op_bot_0')
// (11, 10, 'sp4_r_v_b_20')
// (11, 11, 'sp4_r_v_b_9')
// (12, 5, 'sp4_v_t_36')
// (12, 6, 'sp4_v_b_36')
// (12, 7, 'sp4_h_l_38')
// (12, 7, 'sp4_v_b_25')
// (12, 7, 'sp4_v_t_44')
// (12, 8, 'neigh_op_tnl_0')
// (12, 8, 'sp4_v_b_12')
// (12, 8, 'sp4_v_b_44')
// (12, 9, 'neigh_op_lft_0')
// (12, 9, 'sp4_v_b_1')
// (12, 9, 'sp4_v_b_33')
// (12, 10, 'neigh_op_bnl_0')
// (12, 10, 'sp4_v_b_20')
// (12, 11, 'sp4_v_b_9')

wire n493;
// (8, 7, 'sp4_h_r_4')
// (9, 7, 'local_g0_1')
// (9, 7, 'lutff_0/in_1')
// (9, 7, 'sp4_h_r_17')
// (10, 5, 'neigh_op_tnr_0')
// (10, 6, 'neigh_op_rgt_0')
// (10, 7, 'neigh_op_bnr_0')
// (10, 7, 'sp4_h_r_28')
// (11, 4, 'sp4_r_v_b_41')
// (11, 5, 'neigh_op_top_0')
// (11, 5, 'sp4_r_v_b_28')
// (11, 6, 'lutff_0/out')
// (11, 6, 'sp4_r_v_b_17')
// (11, 7, 'neigh_op_bot_0')
// (11, 7, 'sp4_h_r_41')
// (11, 7, 'sp4_r_v_b_4')
// (12, 3, 'sp4_v_t_41')
// (12, 4, 'sp4_v_b_41')
// (12, 5, 'neigh_op_tnl_0')
// (12, 5, 'sp4_v_b_28')
// (12, 6, 'neigh_op_lft_0')
// (12, 6, 'sp4_v_b_17')
// (12, 7, 'neigh_op_bnl_0')
// (12, 7, 'sp4_h_l_41')
// (12, 7, 'sp4_v_b_4')

reg n494 = 0;
// (8, 7, 'sp4_h_r_7')
// (9, 7, 'local_g0_2')
// (9, 7, 'lutff_4/in_0')
// (9, 7, 'sp4_h_r_18')
// (10, 6, 'neigh_op_tnr_5')
// (10, 7, 'neigh_op_rgt_5')
// (10, 7, 'sp4_h_r_31')
// (10, 8, 'neigh_op_bnr_5')
// (11, 6, 'neigh_op_top_5')
// (11, 7, 'lutff_5/out')
// (11, 7, 'sp4_h_r_42')
// (11, 8, 'neigh_op_bot_5')
// (12, 6, 'neigh_op_tnl_5')
// (12, 7, 'neigh_op_lft_5')
// (12, 7, 'sp4_h_l_42')
// (12, 8, 'neigh_op_bnl_5')

reg n495 = 0;
// (8, 7, 'sp4_h_r_9')
// (9, 7, 'local_g1_4')
// (9, 7, 'lutff_7/in_0')
// (9, 7, 'sp4_h_r_20')
// (10, 6, 'neigh_op_tnr_6')
// (10, 7, 'neigh_op_rgt_6')
// (10, 7, 'sp4_h_r_33')
// (10, 8, 'neigh_op_bnr_6')
// (11, 6, 'neigh_op_top_6')
// (11, 7, 'lutff_6/out')
// (11, 7, 'sp4_h_r_44')
// (11, 8, 'neigh_op_bot_6')
// (12, 6, 'neigh_op_tnl_6')
// (12, 7, 'neigh_op_lft_6')
// (12, 7, 'sp4_h_l_44')
// (12, 8, 'neigh_op_bnl_6')

wire n496;
// (8, 7, 'sp4_r_v_b_40')
// (8, 8, 'neigh_op_tnr_0')
// (8, 8, 'sp4_r_v_b_29')
// (8, 9, 'neigh_op_rgt_0')
// (8, 9, 'sp4_r_v_b_16')
// (8, 10, 'local_g1_0')
// (8, 10, 'local_g1_5')
// (8, 10, 'lutff_1/in_2')
// (8, 10, 'lutff_3/in_3')
// (8, 10, 'neigh_op_bnr_0')
// (8, 10, 'sp4_r_v_b_5')
// (9, 6, 'sp4_v_t_40')
// (9, 7, 'sp4_v_b_40')
// (9, 8, 'neigh_op_top_0')
// (9, 8, 'sp4_v_b_29')
// (9, 9, 'lutff_0/out')
// (9, 9, 'sp4_v_b_16')
// (9, 10, 'local_g1_0')
// (9, 10, 'lutff_4/in_3')
// (9, 10, 'neigh_op_bot_0')
// (9, 10, 'sp4_v_b_5')
// (10, 8, 'neigh_op_tnl_0')
// (10, 9, 'neigh_op_lft_0')
// (10, 10, 'neigh_op_bnl_0')

wire n497;
// (8, 7, 'sp4_r_v_b_42')
// (8, 8, 'neigh_op_tnr_1')
// (8, 8, 'sp4_r_v_b_31')
// (8, 9, 'neigh_op_rgt_1')
// (8, 9, 'sp4_r_v_b_18')
// (8, 10, 'local_g1_1')
// (8, 10, 'lutff_6/in_2')
// (8, 10, 'neigh_op_bnr_1')
// (8, 10, 'sp4_r_v_b_7')
// (8, 11, 'local_g3_2')
// (8, 11, 'lutff_3/in_2')
// (8, 11, 'sp4_r_v_b_42')
// (8, 12, 'sp4_r_v_b_31')
// (8, 13, 'sp4_r_v_b_18')
// (8, 14, 'sp4_r_v_b_7')
// (9, 6, 'sp4_v_t_42')
// (9, 7, 'sp4_v_b_42')
// (9, 8, 'neigh_op_top_1')
// (9, 8, 'sp4_v_b_31')
// (9, 9, 'lutff_1/out')
// (9, 9, 'sp4_v_b_18')
// (9, 10, 'local_g0_7')
// (9, 10, 'lutff_0/in_1')
// (9, 10, 'neigh_op_bot_1')
// (9, 10, 'sp4_v_b_7')
// (9, 10, 'sp4_v_t_42')
// (9, 11, 'local_g2_2')
// (9, 11, 'local_g3_2')
// (9, 11, 'lutff_2/in_2')
// (9, 11, 'lutff_6/in_1')
// (9, 11, 'sp4_v_b_42')
// (9, 12, 'sp4_v_b_31')
// (9, 13, 'sp4_v_b_18')
// (9, 14, 'sp4_v_b_7')
// (10, 8, 'neigh_op_tnl_1')
// (10, 9, 'neigh_op_lft_1')
// (10, 10, 'neigh_op_bnl_1')

wire n498;
// (8, 8, 'neigh_op_tnr_4')
// (8, 9, 'neigh_op_rgt_4')
// (8, 10, 'local_g0_4')
// (8, 10, 'local_g1_4')
// (8, 10, 'lutff_4/in_2')
// (8, 10, 'lutff_6/in_1')
// (8, 10, 'lutff_7/in_1')
// (8, 10, 'neigh_op_bnr_4')
// (9, 8, 'neigh_op_top_4')
// (9, 9, 'lutff_4/out')
// (9, 10, 'local_g1_4')
// (9, 10, 'lutff_2/in_3')
// (9, 10, 'neigh_op_bot_4')
// (10, 8, 'neigh_op_tnl_4')
// (10, 9, 'neigh_op_lft_4')
// (10, 10, 'neigh_op_bnl_4')

wire n499;
// (8, 8, 'neigh_op_tnr_5')
// (8, 9, 'neigh_op_rgt_5')
// (8, 10, 'neigh_op_bnr_5')
// (9, 8, 'neigh_op_top_5')
// (9, 9, 'local_g0_5')
// (9, 9, 'local_g1_5')
// (9, 9, 'lutff_1/in_3')
// (9, 9, 'lutff_4/in_3')
// (9, 9, 'lutff_5/out')
// (9, 10, 'neigh_op_bot_5')
// (10, 8, 'neigh_op_tnl_5')
// (10, 9, 'neigh_op_lft_5')
// (10, 10, 'neigh_op_bnl_5')

reg n500 = 0;
// (8, 8, 'neigh_op_tnr_6')
// (8, 9, 'neigh_op_rgt_6')
// (8, 10, 'neigh_op_bnr_6')
// (9, 8, 'local_g0_6')
// (9, 8, 'lutff_0/in_0')
// (9, 8, 'neigh_op_top_6')
// (9, 9, 'lutff_6/out')
// (9, 10, 'neigh_op_bot_6')
// (10, 8, 'neigh_op_tnl_6')
// (10, 9, 'neigh_op_lft_6')
// (10, 10, 'neigh_op_bnl_6')

wire n501;
// (8, 8, 'sp4_r_v_b_36')
// (8, 9, 'neigh_op_tnr_6')
// (8, 9, 'sp4_r_v_b_25')
// (8, 10, 'neigh_op_rgt_6')
// (8, 10, 'sp4_r_v_b_12')
// (8, 11, 'neigh_op_bnr_6')
// (8, 11, 'sp4_r_v_b_1')
// (9, 7, 'sp4_v_t_36')
// (9, 8, 'sp4_v_b_36')
// (9, 9, 'neigh_op_top_6')
// (9, 9, 'sp4_v_b_25')
// (9, 10, 'lutff_6/out')
// (9, 10, 'sp4_v_b_12')
// (9, 11, 'local_g0_1')
// (9, 11, 'local_g0_6')
// (9, 11, 'lutff_1/in_3')
// (9, 11, 'lutff_4/in_1')
// (9, 11, 'neigh_op_bot_6')
// (9, 11, 'sp4_v_b_1')
// (10, 9, 'neigh_op_tnl_6')
// (10, 10, 'neigh_op_lft_6')
// (10, 11, 'neigh_op_bnl_6')

wire n502;
// (8, 9, 'neigh_op_tnr_0')
// (8, 9, 'sp4_r_v_b_43')
// (8, 10, 'neigh_op_rgt_0')
// (8, 10, 'sp4_r_v_b_30')
// (8, 11, 'neigh_op_bnr_0')
// (8, 11, 'sp4_r_v_b_19')
// (8, 12, 'sp4_r_v_b_6')
// (9, 6, 'sp12_v_t_23')
// (9, 7, 'sp12_v_b_23')
// (9, 8, 'sp12_v_b_20')
// (9, 8, 'sp4_v_t_43')
// (9, 9, 'neigh_op_top_0')
// (9, 9, 'sp12_v_b_19')
// (9, 9, 'sp4_v_b_43')
// (9, 10, 'lutff_0/out')
// (9, 10, 'sp12_v_b_16')
// (9, 10, 'sp4_v_b_30')
// (9, 11, 'local_g1_3')
// (9, 11, 'lutff_5/in_3')
// (9, 11, 'neigh_op_bot_0')
// (9, 11, 'sp12_v_b_15')
// (9, 11, 'sp4_v_b_19')
// (9, 12, 'sp12_v_b_12')
// (9, 12, 'sp4_v_b_6')
// (9, 13, 'sp12_v_b_11')
// (9, 14, 'sp12_v_b_8')
// (9, 15, 'sp12_v_b_7')
// (9, 16, 'sp12_v_b_4')
// (9, 17, 'span12_vert_3')
// (10, 9, 'neigh_op_tnl_0')
// (10, 10, 'neigh_op_lft_0')
// (10, 11, 'neigh_op_bnl_0')

wire n503;
// (8, 9, 'neigh_op_tnr_1')
// (8, 10, 'neigh_op_rgt_1')
// (8, 11, 'neigh_op_bnr_1')
// (9, 9, 'neigh_op_top_1')
// (9, 10, 'local_g0_1')
// (9, 10, 'local_g1_1')
// (9, 10, 'lutff_1/out')
// (9, 10, 'lutff_2/in_2')
// (9, 10, 'lutff_6/in_1')
// (9, 11, 'neigh_op_bot_1')
// (10, 9, 'neigh_op_tnl_1')
// (10, 10, 'neigh_op_lft_1')
// (10, 11, 'neigh_op_bnl_1')

wire n504;
// (8, 9, 'neigh_op_tnr_2')
// (8, 10, 'neigh_op_rgt_2')
// (8, 11, 'neigh_op_bnr_2')
// (9, 8, 'sp4_r_v_b_45')
// (9, 9, 'neigh_op_top_2')
// (9, 9, 'sp4_r_v_b_32')
// (9, 10, 'lutff_2/out')
// (9, 10, 'sp4_r_v_b_21')
// (9, 10, 'sp4_r_v_b_37')
// (9, 11, 'local_g1_0')
// (9, 11, 'local_g2_0')
// (9, 11, 'lutff_4/in_2')
// (9, 11, 'lutff_7/in_2')
// (9, 11, 'neigh_op_bot_2')
// (9, 11, 'sp4_r_v_b_24')
// (9, 11, 'sp4_r_v_b_8')
// (9, 12, 'sp4_r_v_b_13')
// (9, 13, 'sp4_r_v_b_0')
// (10, 7, 'sp4_v_t_45')
// (10, 8, 'sp4_v_b_45')
// (10, 9, 'neigh_op_tnl_2')
// (10, 9, 'sp4_v_b_32')
// (10, 9, 'sp4_v_t_37')
// (10, 10, 'neigh_op_lft_2')
// (10, 10, 'sp4_v_b_21')
// (10, 10, 'sp4_v_b_37')
// (10, 11, 'neigh_op_bnl_2')
// (10, 11, 'sp4_v_b_24')
// (10, 11, 'sp4_v_b_8')
// (10, 12, 'sp4_v_b_13')
// (10, 13, 'sp4_v_b_0')

wire n505;
// (8, 9, 'neigh_op_tnr_4')
// (8, 10, 'neigh_op_rgt_4')
// (8, 11, 'neigh_op_bnr_4')
// (9, 9, 'neigh_op_top_4')
// (9, 10, 'lutff_4/out')
// (9, 11, 'local_g1_4')
// (9, 11, 'lutff_6/in_3')
// (9, 11, 'neigh_op_bot_4')
// (10, 9, 'neigh_op_tnl_4')
// (10, 10, 'neigh_op_lft_4')
// (10, 11, 'neigh_op_bnl_4')

wire n506;
// (8, 9, 'neigh_op_tnr_5')
// (8, 10, 'neigh_op_rgt_5')
// (8, 11, 'local_g1_5')
// (8, 11, 'lutff_0/in_2')
// (8, 11, 'lutff_4/in_2')
// (8, 11, 'neigh_op_bnr_5')
// (9, 9, 'neigh_op_top_5')
// (9, 10, 'local_g0_5')
// (9, 10, 'lutff_2/in_1')
// (9, 10, 'lutff_5/out')
// (9, 11, 'local_g0_5')
// (9, 11, 'local_g1_5')
// (9, 11, 'lutff_2/in_1')
// (9, 11, 'lutff_6/in_0')
// (9, 11, 'neigh_op_bot_5')
// (10, 9, 'neigh_op_tnl_5')
// (10, 10, 'neigh_op_lft_5')
// (10, 11, 'neigh_op_bnl_5')

wire n507;
// (8, 9, 'neigh_op_tnr_7')
// (8, 10, 'neigh_op_rgt_7')
// (8, 11, 'neigh_op_bnr_7')
// (9, 5, 'sp12_v_t_22')
// (9, 6, 'sp12_v_b_22')
// (9, 7, 'sp12_v_b_21')
// (9, 8, 'sp12_v_b_18')
// (9, 9, 'neigh_op_top_7')
// (9, 9, 'sp12_v_b_17')
// (9, 10, 'lutff_7/out')
// (9, 10, 'sp12_v_b_14')
// (9, 11, 'local_g2_5')
// (9, 11, 'lutff_0/in_3')
// (9, 11, 'neigh_op_bot_7')
// (9, 11, 'sp12_v_b_13')
// (9, 12, 'sp12_v_b_10')
// (9, 13, 'sp12_v_b_9')
// (9, 14, 'sp12_v_b_6')
// (9, 15, 'sp12_v_b_5')
// (9, 16, 'sp12_v_b_2')
// (9, 17, 'span12_vert_1')
// (10, 9, 'neigh_op_tnl_7')
// (10, 10, 'neigh_op_lft_7')
// (10, 11, 'neigh_op_bnl_7')

wire n508;
// (8, 10, 'neigh_op_tnr_0')
// (8, 11, 'neigh_op_rgt_0')
// (8, 12, 'neigh_op_bnr_0')
// (9, 10, 'neigh_op_top_0')
// (9, 11, 'local_g0_0')
// (9, 11, 'lutff_0/out')
// (9, 11, 'lutff_1/in_1')
// (9, 12, 'neigh_op_bot_0')
// (10, 10, 'neigh_op_tnl_0')
// (10, 11, 'neigh_op_lft_0')
// (10, 12, 'neigh_op_bnl_0')

wire n509;
// (8, 10, 'neigh_op_tnr_2')
// (8, 11, 'neigh_op_rgt_2')
// (8, 12, 'neigh_op_bnr_2')
// (9, 10, 'neigh_op_top_2')
// (9, 11, 'local_g0_2')
// (9, 11, 'local_g1_2')
// (9, 11, 'lutff_1/in_2')
// (9, 11, 'lutff_2/out')
// (9, 11, 'lutff_5/in_1')
// (9, 11, 'lutff_7/in_1')
// (9, 12, 'neigh_op_bot_2')
// (10, 10, 'neigh_op_tnl_2')
// (10, 11, 'neigh_op_lft_2')
// (10, 12, 'neigh_op_bnl_2')

wire n510;
// (8, 10, 'neigh_op_tnr_3')
// (8, 11, 'neigh_op_rgt_3')
// (8, 12, 'neigh_op_bnr_3')
// (9, 10, 'neigh_op_top_3')
// (9, 11, 'local_g0_3')
// (9, 11, 'lutff_3/out')
// (9, 11, 'lutff_5/in_2')
// (9, 12, 'neigh_op_bot_3')
// (10, 10, 'neigh_op_tnl_3')
// (10, 11, 'neigh_op_lft_3')
// (10, 12, 'neigh_op_bnl_3')

wire n511;
// (8, 10, 'neigh_op_tnr_6')
// (8, 11, 'neigh_op_rgt_6')
// (8, 12, 'neigh_op_bnr_6')
// (9, 10, 'neigh_op_top_6')
// (9, 11, 'local_g1_6')
// (9, 11, 'lutff_4/in_3')
// (9, 11, 'lutff_6/out')
// (9, 12, 'neigh_op_bot_6')
// (10, 10, 'neigh_op_tnl_6')
// (10, 11, 'neigh_op_lft_6')
// (10, 12, 'neigh_op_bnl_6')

wire n512;
// (8, 12, 'neigh_op_tnr_0')
// (8, 13, 'neigh_op_rgt_0')
// (8, 14, 'neigh_op_bnr_0')
// (9, 12, 'neigh_op_top_0')
// (9, 13, 'local_g1_0')
// (9, 13, 'lutff_0/out')
// (9, 13, 'lutff_2/in_3')
// (9, 14, 'neigh_op_bot_0')
// (10, 12, 'neigh_op_tnl_0')
// (10, 13, 'neigh_op_lft_0')
// (10, 14, 'neigh_op_bnl_0')

wire n513;
// (8, 12, 'neigh_op_tnr_2')
// (8, 13, 'local_g2_2')
// (8, 13, 'lutff_4/in_2')
// (8, 13, 'neigh_op_rgt_2')
// (8, 14, 'neigh_op_bnr_2')
// (9, 12, 'neigh_op_top_2')
// (9, 13, 'lutff_2/out')
// (9, 14, 'neigh_op_bot_2')
// (10, 12, 'neigh_op_tnl_2')
// (10, 13, 'neigh_op_lft_2')
// (10, 14, 'neigh_op_bnl_2')

reg n514 = 0;
// (10, 3, 'neigh_op_tnr_3')
// (10, 4, 'neigh_op_rgt_3')
// (10, 5, 'neigh_op_bnr_3')
// (11, 3, 'neigh_op_top_3')
// (11, 4, 'lutff_3/out')
// (11, 5, 'local_g0_3')
// (11, 5, 'lutff_5/in_0')
// (11, 5, 'neigh_op_bot_3')
// (12, 3, 'neigh_op_tnl_3')
// (12, 4, 'neigh_op_lft_3')
// (12, 5, 'neigh_op_bnl_3')

reg n515 = 0;
// (10, 4, 'neigh_op_tnr_5')
// (10, 5, 'neigh_op_rgt_5')
// (10, 6, 'neigh_op_bnr_5')
// (11, 4, 'neigh_op_top_5')
// (11, 5, 'local_g1_5')
// (11, 5, 'lutff_5/out')
// (11, 5, 'lutff_6/in_0')
// (11, 6, 'neigh_op_bot_5')
// (12, 4, 'neigh_op_tnl_5')
// (12, 5, 'neigh_op_lft_5')
// (12, 6, 'neigh_op_bnl_5')

reg n516 = 0;
// (10, 5, 'neigh_op_tnr_3')
// (10, 6, 'neigh_op_rgt_3')
// (10, 7, 'neigh_op_bnr_3')
// (11, 5, 'neigh_op_top_3')
// (11, 6, 'local_g1_3')
// (11, 6, 'lutff_3/out')
// (11, 6, 'lutff_4/in_0')
// (11, 7, 'neigh_op_bot_3')
// (12, 5, 'neigh_op_tnl_3')
// (12, 6, 'neigh_op_lft_3')
// (12, 7, 'neigh_op_bnl_3')

reg n517 = 0;
// (10, 5, 'neigh_op_tnr_5')
// (10, 6, 'neigh_op_rgt_5')
// (10, 7, 'neigh_op_bnr_5')
// (11, 5, 'neigh_op_top_5')
// (11, 6, 'local_g0_5')
// (11, 6, 'lutff_3/in_0')
// (11, 6, 'lutff_5/out')
// (11, 7, 'neigh_op_bot_5')
// (12, 5, 'neigh_op_tnl_5')
// (12, 6, 'neigh_op_lft_5')
// (12, 7, 'neigh_op_bnl_5')

reg n518 = 0;
// (10, 5, 'neigh_op_tnr_6')
// (10, 6, 'neigh_op_rgt_6')
// (10, 7, 'neigh_op_bnr_6')
// (11, 5, 'neigh_op_top_6')
// (11, 6, 'local_g1_6')
// (11, 6, 'lutff_6/out')
// (11, 6, 'lutff_7/in_0')
// (11, 7, 'neigh_op_bot_6')
// (12, 5, 'neigh_op_tnl_6')
// (12, 6, 'neigh_op_lft_6')
// (12, 7, 'neigh_op_bnl_6')

reg n519 = 0;
// (10, 6, 'neigh_op_tnr_2')
// (10, 7, 'neigh_op_rgt_2')
// (10, 8, 'neigh_op_bnr_2')
// (11, 6, 'neigh_op_top_2')
// (11, 7, 'local_g1_2')
// (11, 7, 'lutff_2/out')
// (11, 7, 'lutff_5/in_0')
// (11, 8, 'neigh_op_bot_2')
// (12, 6, 'neigh_op_tnl_2')
// (12, 7, 'neigh_op_lft_2')
// (12, 8, 'neigh_op_bnl_2')

reg n520 = 0;
// (10, 6, 'neigh_op_tnr_4')
// (10, 7, 'neigh_op_rgt_4')
// (10, 8, 'neigh_op_bnr_4')
// (11, 6, 'neigh_op_top_4')
// (11, 7, 'local_g0_4')
// (11, 7, 'lutff_4/out')
// (11, 7, 'lutff_6/in_0')
// (11, 8, 'neigh_op_bot_4')
// (12, 6, 'neigh_op_tnl_4')
// (12, 7, 'neigh_op_lft_4')
// (12, 8, 'neigh_op_bnl_4')

reg n521 = 0;
// (10, 6, 'neigh_op_tnr_7')
// (10, 7, 'neigh_op_rgt_7')
// (10, 8, 'neigh_op_bnr_7')
// (11, 6, 'neigh_op_top_7')
// (11, 7, 'local_g0_7')
// (11, 7, 'lutff_0/in_1')
// (11, 7, 'lutff_7/out')
// (11, 8, 'neigh_op_bot_7')
// (12, 6, 'neigh_op_tnl_7')
// (12, 7, 'neigh_op_lft_7')
// (12, 8, 'neigh_op_bnl_7')

reg n522 = 0;
// (10, 7, 'neigh_op_tnr_3')
// (10, 8, 'neigh_op_rgt_3')
// (10, 9, 'neigh_op_bnr_3')
// (11, 6, 'sp4_r_v_b_47')
// (11, 7, 'local_g2_2')
// (11, 7, 'lutff_7/in_1')
// (11, 7, 'neigh_op_top_3')
// (11, 7, 'sp4_r_v_b_34')
// (11, 8, 'lutff_3/out')
// (11, 8, 'sp4_r_v_b_23')
// (11, 9, 'neigh_op_bot_3')
// (11, 9, 'sp4_r_v_b_10')
// (12, 5, 'sp4_v_t_47')
// (12, 6, 'sp4_v_b_47')
// (12, 7, 'neigh_op_tnl_3')
// (12, 7, 'sp4_v_b_34')
// (12, 8, 'neigh_op_lft_3')
// (12, 8, 'sp4_v_b_23')
// (12, 9, 'neigh_op_bnl_3')
// (12, 9, 'sp4_v_b_10')

reg n523 = 0;
// (10, 8, 'neigh_op_tnr_1')
// (10, 9, 'neigh_op_rgt_1')
// (10, 10, 'neigh_op_bnr_1')
// (11, 8, 'neigh_op_top_1')
// (11, 9, 'local_g0_1')
// (11, 9, 'lutff_1/out')
// (11, 9, 'lutff_2/in_1')
// (11, 10, 'neigh_op_bot_1')
// (12, 8, 'neigh_op_tnl_1')
// (12, 9, 'neigh_op_lft_1')
// (12, 10, 'neigh_op_bnl_1')

reg n524 = 0;
// (10, 8, 'neigh_op_tnr_2')
// (10, 9, 'neigh_op_rgt_2')
// (10, 10, 'neigh_op_bnr_2')
// (11, 8, 'neigh_op_top_2')
// (11, 9, 'local_g1_2')
// (11, 9, 'lutff_0/in_1')
// (11, 9, 'lutff_2/out')
// (11, 10, 'neigh_op_bot_2')
// (12, 8, 'neigh_op_tnl_2')
// (12, 9, 'neigh_op_lft_2')
// (12, 10, 'neigh_op_bnl_2')

reg n525 = 0;
// (10, 8, 'neigh_op_tnr_4')
// (10, 9, 'neigh_op_rgt_4')
// (10, 10, 'neigh_op_bnr_4')
// (11, 8, 'neigh_op_top_4')
// (11, 9, 'local_g0_4')
// (11, 9, 'lutff_0/in_0')
// (11, 9, 'lutff_4/out')
// (11, 9, 'lutff_7/in_1')
// (11, 10, 'neigh_op_bot_4')
// (12, 8, 'neigh_op_tnl_4')
// (12, 9, 'neigh_op_lft_4')
// (12, 10, 'neigh_op_bnl_4')

reg n526 = 0;
// (10, 8, 'neigh_op_tnr_5')
// (10, 9, 'neigh_op_rgt_5')
// (10, 10, 'neigh_op_bnr_5')
// (11, 8, 'neigh_op_top_5')
// (11, 9, 'local_g0_5')
// (11, 9, 'local_g3_5')
// (11, 9, 'lutff_2/in_2')
// (11, 9, 'lutff_4/in_1')
// (11, 9, 'lutff_5/out')
// (11, 10, 'neigh_op_bot_5')
// (12, 8, 'neigh_op_tnl_5')
// (12, 9, 'neigh_op_lft_5')
// (12, 10, 'neigh_op_bnl_5')

reg n527 = 0;
// (10, 8, 'neigh_op_tnr_6')
// (10, 9, 'neigh_op_rgt_6')
// (10, 10, 'neigh_op_bnr_6')
// (11, 8, 'neigh_op_top_6')
// (11, 9, 'local_g0_6')
// (11, 9, 'local_g1_6')
// (11, 9, 'lutff_1/in_2')
// (11, 9, 'lutff_5/in_1')
// (11, 9, 'lutff_6/out')
// (11, 10, 'neigh_op_bot_6')
// (12, 8, 'neigh_op_tnl_6')
// (12, 9, 'neigh_op_lft_6')
// (12, 10, 'neigh_op_bnl_6')

reg n528 = 0;
// (10, 8, 'neigh_op_tnr_7')
// (10, 9, 'neigh_op_rgt_7')
// (10, 10, 'neigh_op_bnr_7')
// (11, 8, 'neigh_op_top_7')
// (11, 9, 'local_g0_7')
// (11, 9, 'lutff_6/in_1')
// (11, 9, 'lutff_7/out')
// (11, 10, 'neigh_op_bot_7')
// (12, 8, 'neigh_op_tnl_7')
// (12, 9, 'local_g1_7')
// (12, 9, 'lutff_6/in_0')
// (12, 9, 'neigh_op_lft_7')
// (12, 10, 'neigh_op_bnl_7')

wire n529;
// (10, 10, 'neigh_op_tnr_0')
// (10, 11, 'neigh_op_rgt_0')
// (10, 12, 'neigh_op_bnr_0')
// (11, 10, 'local_g1_0')
// (11, 10, 'lutff_4/in_3')
// (11, 10, 'neigh_op_top_0')
// (11, 11, 'local_g1_0')
// (11, 11, 'lutff_0/out')
// (11, 11, 'lutff_5/in_0')
// (11, 12, 'neigh_op_bot_0')
// (12, 10, 'neigh_op_tnl_0')
// (12, 11, 'neigh_op_lft_0')
// (12, 12, 'neigh_op_bnl_0')

reg n530 = 0;
// (10, 10, 'sp4_r_v_b_41')
// (10, 11, 'sp4_r_v_b_28')
// (10, 12, 'neigh_op_tnr_2')
// (10, 12, 'sp4_r_v_b_17')
// (10, 13, 'neigh_op_rgt_2')
// (10, 13, 'sp4_r_v_b_4')
// (10, 14, 'neigh_op_bnr_2')
// (11, 9, 'sp4_v_t_41')
// (11, 10, 'sp4_v_b_41')
// (11, 11, 'local_g2_4')
// (11, 11, 'lutff_4/in_2')
// (11, 11, 'sp4_v_b_28')
// (11, 12, 'local_g1_2')
// (11, 12, 'lutff_4/in_1')
// (11, 12, 'neigh_op_top_2')
// (11, 12, 'sp4_v_b_17')
// (11, 13, 'local_g0_2')
// (11, 13, 'lutff_2/in_2')
// (11, 13, 'lutff_2/out')
// (11, 13, 'sp4_v_b_4')
// (11, 14, 'neigh_op_bot_2')
// (12, 12, 'neigh_op_tnl_2')
// (12, 13, 'neigh_op_lft_2')
// (12, 14, 'neigh_op_bnl_2')

wire n531;
// (10, 11, 'neigh_op_tnr_1')
// (10, 12, 'neigh_op_rgt_1')
// (10, 13, 'neigh_op_bnr_1')
// (11, 11, 'neigh_op_top_1')
// (11, 12, 'local_g0_1')
// (11, 12, 'lutff_1/out')
// (11, 12, 'lutff_3/in_2')
// (11, 13, 'neigh_op_bot_1')
// (12, 11, 'neigh_op_tnl_1')
// (12, 12, 'neigh_op_lft_1')
// (12, 13, 'neigh_op_bnl_1')

wire n532;
// (10, 11, 'neigh_op_tnr_3')
// (10, 12, 'neigh_op_rgt_3')
// (10, 13, 'neigh_op_bnr_3')
// (11, 11, 'neigh_op_top_3')
// (11, 12, 'lutff_3/out')
// (11, 13, 'neigh_op_bot_3')
// (12, 11, 'neigh_op_tnl_3')
// (12, 12, 'local_g1_3')
// (12, 12, 'lutff_global/cen')
// (12, 12, 'neigh_op_lft_3')
// (12, 13, 'neigh_op_bnl_3')

wire n533;
// (10, 11, 'neigh_op_tnr_4')
// (10, 12, 'neigh_op_rgt_4')
// (10, 13, 'neigh_op_bnr_4')
// (11, 11, 'neigh_op_top_4')
// (11, 12, 'local_g0_4')
// (11, 12, 'lutff_3/in_1')
// (11, 12, 'lutff_4/out')
// (11, 13, 'neigh_op_bot_4')
// (12, 11, 'neigh_op_tnl_4')
// (12, 12, 'neigh_op_lft_4')
// (12, 13, 'neigh_op_bnl_4')

reg n534 = 0;
// (10, 12, 'neigh_op_tnr_3')
// (10, 13, 'neigh_op_rgt_3')
// (10, 14, 'neigh_op_bnr_3')
// (11, 10, 'sp4_r_v_b_42')
// (11, 11, 'local_g0_7')
// (11, 11, 'local_g1_7')
// (11, 11, 'lutff_4/in_1')
// (11, 11, 'lutff_7/in_1')
// (11, 11, 'sp4_r_v_b_31')
// (11, 12, 'local_g0_3')
// (11, 12, 'lutff_4/in_3')
// (11, 12, 'neigh_op_top_3')
// (11, 12, 'sp4_r_v_b_18')
// (11, 13, 'local_g0_3')
// (11, 13, 'lutff_3/in_2')
// (11, 13, 'lutff_3/out')
// (11, 13, 'sp4_r_v_b_7')
// (11, 14, 'neigh_op_bot_3')
// (12, 9, 'sp4_v_t_42')
// (12, 10, 'sp4_v_b_42')
// (12, 11, 'sp4_v_b_31')
// (12, 12, 'neigh_op_tnl_3')
// (12, 12, 'sp4_v_b_18')
// (12, 13, 'neigh_op_lft_3')
// (12, 13, 'sp4_v_b_7')
// (12, 14, 'neigh_op_bnl_3')

reg n535 = 0;
// (11, 6, 'neigh_op_tnr_1')
// (11, 7, 'neigh_op_rgt_1')
// (11, 8, 'neigh_op_bnr_1')
// (12, 6, 'neigh_op_top_1')
// (12, 7, 'local_g1_1')
// (12, 7, 'lutff_1/out')
// (12, 7, 'lutff_6/in_0')
// (12, 8, 'neigh_op_bot_1')
// (13, 6, 'logic_op_tnl_1')
// (13, 7, 'logic_op_lft_1')
// (13, 8, 'logic_op_bnl_1')

reg n536 = 0;
// (11, 6, 'neigh_op_tnr_6')
// (11, 7, 'neigh_op_rgt_6')
// (11, 8, 'neigh_op_bnr_6')
// (12, 6, 'neigh_op_top_6')
// (12, 7, 'local_g1_6')
// (12, 7, 'lutff_3/in_0')
// (12, 7, 'lutff_6/out')
// (12, 8, 'neigh_op_bot_6')
// (13, 6, 'logic_op_tnl_6')
// (13, 7, 'logic_op_lft_6')
// (13, 8, 'logic_op_bnl_6')

reg n537 = 0;
// (11, 8, 'neigh_op_tnr_6')
// (11, 9, 'local_g2_6')
// (11, 9, 'lutff_1/in_1')
// (11, 9, 'neigh_op_rgt_6')
// (11, 10, 'neigh_op_bnr_6')
// (12, 8, 'neigh_op_top_6')
// (12, 9, 'lutff_6/out')
// (12, 10, 'neigh_op_bot_6')
// (13, 8, 'logic_op_tnl_6')
// (13, 9, 'logic_op_lft_6')
// (13, 10, 'logic_op_bnl_6')

reg d_vld = 0;
// (11, 10, 'sp4_r_v_b_40')
// (11, 11, 'neigh_op_tnr_0')
// (11, 11, 'sp4_r_v_b_29')
// (11, 12, 'neigh_op_rgt_0')
// (11, 12, 'sp4_r_v_b_16')
// (11, 13, 'neigh_op_bnr_0')
// (11, 13, 'sp4_r_v_b_5')
// (12, 9, 'sp4_h_r_5')
// (12, 9, 'sp4_v_t_40')
// (12, 10, 'sp4_v_b_40')
// (12, 11, 'neigh_op_top_0')
// (12, 11, 'sp4_v_b_29')
// (12, 12, 'lutff_0/out')
// (12, 12, 'sp4_v_b_16')
// (12, 13, 'neigh_op_bot_0')
// (12, 13, 'sp4_v_b_5')
// (13, 9, 'io_1/D_OUT_0')
// (13, 9, 'io_1/PAD')
// (13, 9, 'local_g0_5')
// (13, 9, 'span4_horz_5')
// (13, 11, 'logic_op_tnl_0')
// (13, 12, 'logic_op_lft_0')
// (13, 13, 'logic_op_bnl_0')

wire n539;
// (11, 13, 'lutff_1/cout')
// (11, 13, 'lutff_2/in_3')

wire n540;
// (11, 13, 'lutff_2/cout')
// (11, 13, 'lutff_3/in_3')

wire n541;
// (11, 13, 'lutff_3/cout')
// (11, 13, 'lutff_4/in_3')

wire n542;
// (11, 13, 'lutff_4/cout')
// (11, 13, 'lutff_5/in_3')

wire n543;
// (11, 13, 'lutff_5/cout')
// (11, 13, 'lutff_6/in_3')

wire n544;
// (11, 13, 'lutff_6/cout')
// (11, 13, 'lutff_7/in_3')

wire n545;
// (4, 14, 'lutff_0/cout')

wire n546;
// (11, 13, 'lutff_0/cout')

wire n547;
// (5, 12, 'lutff_6/lout')

wire n548;
// (9, 12, 'lutff_1/lout')

wire n549;
// (5, 4, 'lutff_2/lout')

wire n550;
// (4, 8, 'lutff_5/lout')

wire n551;
// (8, 8, 'lutff_6/lout')

wire n552;
// (7, 4, 'lutff_4/lout')

wire n553;
// (7, 13, 'lutff_0/lout')

wire n554;
// (9, 13, 'lutff_2/lout')

wire n555;
// (5, 5, 'lutff_3/lout')

wire n556;
// (6, 12, 'lutff_1/lout')

wire n557;
// (7, 5, 'lutff_5/lout')

wire n558;
// (4, 12, 'lutff_2/lout')

wire n559;
// (8, 12, 'lutff_3/lout')

wire n560;
// (6, 15, 'lutff_3/lout')

wire n561;
// (5, 9, 'lutff_0/lout')

wire n562;
// (9, 9, 'lutff_4/lout')

wire n563;
// (5, 8, 'lutff_4/lout')

wire n564;
// (7, 8, 'lutff_6/lout')

wire n565;
// (4, 15, 'lutff_3/lout')

wire n566;
// (11, 6, 'lutff_5/lout')

wire n567;
// (8, 11, 'lutff_7/lout')

wire n568;
// (5, 12, 'lutff_1/lout')

wire n569;
// (7, 12, 'lutff_3/lout')

wire n570;
// (4, 8, 'lutff_0/lout')

wire n571;
// (8, 8, 'lutff_1/lout')

wire n572;
// (5, 4, 'lutff_6/lout')

wire n573;
// (7, 13, 'lutff_4/lout')

wire n574;
// (7, 5, 'lutff_0/lout')

wire n575;
// (5, 5, 'lutff_7/lout')

wire n576;
// (9, 5, 'lutff_2/lout')

wire n577;
// (2, 12, 'lutff_4/lout')

wire n578;
// (2, 4, 'lutff_0/lout')

wire n579;
// (4, 12, 'lutff_6/lout')

wire n580;
// (6, 15, 'lutff_7/lout')

wire n581;
// (6, 7, 'lutff_3/lout')

wire n582;
// (7, 8, 'lutff_1/lout')

wire n583;
// (5, 11, 'lutff_4/lout')

wire n584;
// (4, 15, 'lutff_7/lout')

wire n585;
// (7, 11, 'lutff_6/lout')

wire n586;
// (4, 7, 'lutff_3/lout')

wire n587;
// (11, 6, 'lutff_0/lout')

wire n588;
// (8, 11, 'lutff_2/lout')

wire n589;
// (11, 9, 'lutff_5/lout')

wire n590;
// (5, 12, 'lutff_5/lout')

wire n591;
// (7, 12, 'lutff_7/lout')

wire n592;
// (5, 4, 'lutff_1/lout')

wire n593;
// (6, 8, 'lutff_3/lout')

wire n594;
// (4, 8, 'lutff_4/lout')

wire n595;
// (7, 4, 'lutff_3/lout')

wire n596;
// (8, 8, 'lutff_5/lout')

wire n597;
// (6, 3, 'lutff_1/lout')

wire n598;
// (6, 14, 'lutff_1/lout')

wire n599;
// (8, 3, 'lutff_3/lout')

wire n600;
// (6, 6, 'lutff_6/lout')

wire n601;
// (4, 11, 'lutff_5/lout')

wire n602;
// (6, 15, 'lutff_2/lout')

wire n603;
// (8, 7, 'lutff_0/lout')

wire n604;
// (6, 7, 'lutff_7/lout')

wire n605;
// (11, 13, 'lutff_7/lout')

wire n606;
// (5, 8, 'lutff_3/lout')

wire n607;
// (7, 8, 'lutff_5/lout')

wire n608;
// (4, 15, 'lutff_2/lout')

wire n609;
// (9, 8, 'lutff_7/lout')

wire n610;
// (7, 11, 'lutff_1/lout')

wire n611;
// (4, 7, 'lutff_7/lout')

wire n612;
// (6, 11, 'lutff_4/lout')

wire n613;
// (8, 11, 'lutff_6/lout')

wire n614;
// (11, 6, 'lutff_4/lout')

wire n615;
// (11, 9, 'lutff_0/lout')

wire n616;
// (5, 12, 'lutff_0/lout')

wire n617;
// (7, 12, 'lutff_2/lout')

wire n618;
// (5, 4, 'lutff_5/lout')

wire n619;
// (2, 11, 'lutff_2/lout')

wire n620;
// (7, 4, 'lutff_7/lout')

wire n621;
// (6, 3, 'lutff_5/lout')

wire n622;
// (6, 14, 'lutff_5/lout')

wire n623;
// (8, 14, 'lutff_7/lout')

wire n624;
// (6, 6, 'lutff_1/lout')

wire n625;
// (8, 3, 'lutff_7/lout')

wire n626;
// (4, 11, 'lutff_0/lout')

wire n627;
// (5, 7, 'lutff_6/lout')

wire n628;
// (9, 7, 'lutff_1/lout')

wire n629;
// (2, 3, 'lutff_3/lout')

wire n630;
// (4, 14, 'lutff_5/lout')

wire n631;
// (6, 7, 'lutff_2/lout')

wire n632;
// (11, 13, 'lutff_2/lout')

wire n633;
// (5, 8, 'lutff_7/lout')

wire n634;
// (9, 8, 'lutff_2/lout')

wire n635;
// (5, 11, 'lutff_3/lout')

wire n636;
// (2, 7, 'lutff_0/lout')

wire n637;
// (4, 15, 'lutff_6/lout')

wire n638;
// (4, 7, 'lutff_2/lout')

wire n639;
// (8, 11, 'lutff_1/lout')

wire n640;
// (6, 10, 'lutff_3/lout')

wire n641;
// (11, 9, 'lutff_4/lout')

wire n642;
// (8, 10, 'lutff_5/lout')

wire n643;
// (5, 4, 'lutff_0/lout')

wire n644;
// (7, 4, 'lutff_2/lout')

wire n645;
// (9, 11, 'lutff_3/lout')

wire n646;
// (7, 3, 'lutff_6/lout')

wire n647;
// (4, 10, 'lutff_3/lout')

wire n648;
// (6, 3, 'lutff_0/lout')

wire n649;
// (6, 14, 'lutff_0/lout')

wire n650;
// (8, 14, 'lutff_2/lout')

wire n651;
// (8, 3, 'lutff_2/lout')

wire n652;
// (6, 6, 'lutff_5/lout')

wire n653;
// (11, 12, 'lutff_5/lout')

wire n654;
// (9, 4, 'lutff_0/lout')

wire n655;
// (5, 7, 'lutff_1/lout')

wire n656;
// (7, 15, 'lutff_7/lout')

wire n657;
// (4, 11, 'lutff_4/lout')

wire n658;
// (6, 15, 'lutff_1/lout')

wire n659;
// (7, 7, 'lutff_3/lout')

wire n660;
// (4, 3, 'lutff_0/lout')

wire n661;
// (9, 7, 'lutff_5/lout')

wire n662;
// (4, 14, 'lutff_0/out')

wire n663;
// (4, 14, 'lutff_0/lout')

wire n664;
// (4, 14, 'carry_in_mux')

// Carry-In for (4 14)
assign n664 = 1;

wire n665;
// (11, 13, 'lutff_6/lout')

wire n666;
// (12, 12, 'lutff_0/lout')

wire n667;
// (5, 8, 'lutff_2/lout')

wire n668;
// (4, 15, 'lutff_1/lout')

wire n669;
// (4, 4, 'lutff_1/lout')

wire n670;
// (7, 11, 'lutff_0/lout')

wire n671;
// (4, 7, 'lutff_6/lout')

wire n672;
// (11, 6, 'lutff_3/lout')

wire n673;
// (8, 10, 'lutff_0/lout')

wire n674;
// (6, 10, 'lutff_7/lout')

wire n675;
// (6, 13, 'lutff_3/lout')

wire n676;
// (7, 3, 'lutff_1/lout')

wire n677;
// (9, 11, 'lutff_7/lout')

wire n678;
// (9, 3, 'lutff_3/lout')

wire n679;
// (5, 6, 'lutff_4/lout')

wire n680;
// (6, 3, 'lutff_4/lout')

wire n681;
// (6, 14, 'lutff_4/lout')

wire n682;
// (8, 3, 'lutff_6/lout')

wire n683;
// (8, 14, 'lutff_6/lout')

wire n684;
// (5, 15, 'lutff_0/lout')

wire n685;
// (7, 15, 'lutff_2/lout')

wire n686;
// (9, 4, 'lutff_4/lout')

wire n687;
// (5, 7, 'lutff_5/lout')

wire n688;
// (9, 7, 'lutff_0/lout')

wire n689;
// (7, 7, 'lutff_7/lout')

wire n690;
// (4, 3, 'lutff_4/lout')

wire n691;
// (4, 14, 'lutff_4/lout')

wire n692;
// (11, 13, 'lutff_1/out')

wire n693;
// (11, 13, 'lutff_1/lout')

wire n694;
// (11, 5, 'lutff_6/lout')

wire n695;
// (6, 9, 'lutff_1/lout')

wire n696;
// (8, 6, 'lutff_7/lout')

wire n697;
// (7, 14, 'lutff_6/lout')

wire n698;
// (8, 10, 'lutff_4/lout')

wire n699;
// (6, 13, 'lutff_7/lout')

wire n700;
// (6, 2, 'lutff_7/lout')

wire n701;
// (9, 11, 'lutff_2/lout')

wire n702;
// (5, 3, 'lutff_3/lout')

wire n703;
// (4, 10, 'lutff_2/lout')

wire n704;
// (8, 3, 'lutff_1/lout')

wire n705;
// (8, 14, 'lutff_1/lout')

wire n706;
// (6, 6, 'lutff_4/lout')

wire n707;
// (11, 12, 'lutff_4/lout')

wire n708;
// (5, 7, 'lutff_0/lout')

wire n709;
// (7, 15, 'lutff_6/lout')

wire n710;
// (7, 7, 'lutff_2/lout')

wire n711;
// (9, 7, 'lutff_4/lout')

wire n712;
// (5, 10, 'lutff_2/lout')

wire n713;
// (7, 10, 'lutff_4/lout')

wire n714;
// (8, 6, 'lutff_2/lout')

wire n715;
// (9, 10, 'lutff_6/lout')

wire n716;
// (6, 9, 'lutff_5/lout')

wire n717;
// (8, 9, 'lutff_7/lout')

wire n718;
// (7, 14, 'lutff_1/lout')

wire n719;
// (12, 7, 'lutff_6/lout')

wire n720;
// (6, 10, 'lutff_6/lout')

wire n721;
// (6, 13, 'lutff_2/lout')

wire n722;
// (9, 11, 'lutff_6/lout')

wire n723;
// (7, 3, 'lutff_0/lout')

wire n724;
// (5, 3, 'lutff_7/lout')

wire n725;
// (5, 6, 'lutff_3/lout')

wire n726;
// (4, 10, 'lutff_6/lout')

wire n727;
// (8, 13, 'lutff_0/lout')

wire n728;
// (6, 5, 'lutff_3/lout')

wire n729;
// (8, 5, 'lutff_5/lout')

wire n730;
// (5, 10, 'lutff_6/lout')

wire n731;
// (9, 10, 'lutff_1/lout')

wire n732;
// (6, 9, 'lutff_0/lout')

wire n733;
// (8, 6, 'lutff_6/lout')

wire n734;
// (11, 7, 'lutff_5/lout')

wire n735;
// (12, 7, 'lutff_1/lout')

wire n736;
// (6, 10, 'lutff_1/lout')

wire n737;
// (7, 14, 'lutff_5/lout')

wire n738;
// (8, 10, 'lutff_3/lout')

wire n739;
// (6, 13, 'lutff_6/lout')

wire n740;
// (9, 11, 'lutff_1/lout')

wire n741;
// (5, 3, 'lutff_2/lout')

wire n742;
// (7, 3, 'lutff_4/lout')

wire n743;
// (9, 3, 'lutff_6/lout')

wire n744;
// (5, 6, 'lutff_7/lout')

wire n745;
// (7, 6, 'lutff_6/lout')

wire n746;
// (11, 12, 'lutff_3/lout')

wire n747;
// (8, 13, 'lutff_4/lout')

wire n748;
// (8, 5, 'lutff_0/lout')

wire n749;
// (6, 5, 'lutff_7/lout')

wire n750;
// (11, 11, 'lutff_7/lout')

wire n751;
// (5, 10, 'lutff_1/lout')

wire n752;
// (7, 10, 'lutff_3/lout')

wire n753;
// (8, 6, 'lutff_1/lout')

wire n754;
// (9, 10, 'lutff_5/lout')

wire n755;
// (6, 9, 'lutff_4/lout')

wire n756;
// (4, 9, 'lutff_5/lout')

wire n757;
// (8, 9, 'lutff_6/lout')

wire n758;
// (11, 7, 'lutff_0/lout')

wire n759;
// (7, 14, 'lutff_0/lout')

wire n760;
// (11, 8, 'lutff_1/lout')

wire n761;
// (6, 12, 'lutff_5/lout')

wire n762;
// (8, 12, 'lutff_7/lout')

wire n763;
// (7, 6, 'lutff_1/lout')

wire n764;
// (9, 6, 'lutff_3/lout')

wire n765;
// (5, 9, 'lutff_4/lout')

wire n766;
// (4, 13, 'lutff_7/lout')

wire n767;
// (2, 5, 'lutff_1/lout')

wire n768;
// (7, 9, 'lutff_6/lout')

wire n769;
// (6, 5, 'lutff_2/lout')

wire n770;
// (8, 5, 'lutff_4/lout')

wire n771;
// (5, 10, 'lutff_5/lout')

wire n772;
// (9, 10, 'lutff_0/lout')

wire n773;
// (7, 10, 'lutff_7/lout')

wire n774;
// (8, 9, 'lutff_1/lout')

wire n775;
// (11, 7, 'lutff_4/lout')

wire n776;
// (4, 6, 'lutff_3/lout')

wire n777;
// (5, 5, 'lutff_2/lout')

wire n778;
// (6, 12, 'lutff_0/lout')

wire n779;
// (7, 5, 'lutff_4/lout')

wire n780;
// (4, 12, 'lutff_1/lout')

wire n781;
// (8, 12, 'lutff_2/lout')

wire n782;
// (9, 5, 'lutff_6/lout')

wire n783;
// (8, 4, 'lutff_7/lout')

wire n784;
// (7, 6, 'lutff_5/lout')

wire n785;
// (8, 13, 'lutff_3/lout')

wire n786;
// (7, 9, 'lutff_1/lout')

wire n787;
// (9, 6, 'lutff_7/lout')

wire n788;
// (6, 5, 'lutff_6/lout')

wire n789;
// (5, 10, 'lutff_0/lout')

wire n790;
// (7, 10, 'lutff_2/lout')

wire n791;
// (9, 10, 'lutff_4/lout')

wire n792;
// (8, 8, 'lutff_0/lout')

wire n793;
// (2, 8, 'lutff_6/lout')

wire n794;
// (6, 8, 'lutff_7/lout')

wire n795;
// (7, 13, 'lutff_3/lout')

wire n796;
// (9, 13, 'lutff_5/lout')

wire n797;
// (5, 5, 'lutff_6/lout')

wire n798;
// (9, 5, 'lutff_1/lout')

wire n799;
// (6, 12, 'lutff_4/lout')

wire n800;
// (4, 12, 'lutff_5/lout')

wire n801;
// (6, 4, 'lutff_0/lout')

wire n802;
// (8, 12, 'lutff_6/lout')

wire n803;
// (8, 4, 'lutff_2/lout')

wire n804;
// (7, 6, 'lutff_0/lout')

wire n805;
// (9, 6, 'lutff_2/lout')

wire n806;
// (5, 9, 'lutff_3/lout')

wire n807;
// (7, 9, 'lutff_5/lout')

wire n808;
// (6, 5, 'lutff_1/lout')

wire n809;
// (8, 5, 'lutff_3/lout')

wire n810;
// (5, 12, 'lutff_4/lout')

wire n811;
// (7, 1, 'lutff_6/lout')

wire n812;
// (6, 8, 'lutff_2/lout')

wire n813;
// (7, 12, 'lutff_6/lout')

wire n814;
// (4, 8, 'lutff_3/lout')

wire n815;
// (8, 8, 'lutff_4/lout')

wire n816;
// (2, 11, 'lutff_6/lout')

wire n817;
// (9, 13, 'lutff_0/lout')

wire n818;
// (5, 5, 'lutff_1/lout')

wire n819;
// (7, 13, 'lutff_7/lout')

wire n820;
// (8, 12, 'lutff_1/lout')

wire n821;
// (2, 12, 'lutff_7/lout')

wire n822;
// (9, 5, 'lutff_5/lout')

wire n823;
// (6, 4, 'lutff_4/lout')

wire n824;
// (6, 7, 'lutff_6/lout')

wire n825;
// (9, 6, 'lutff_6/lout')

wire n826;
// (7, 9, 'lutff_0/lout')

wire n827;
// (11, 11, 'lutff_5/lout')

wire n828;
// (11, 3, 'lutff_1/lout')

wire n829;
// (6, 11, 'lutff_3/lout')

wire n830;
// (8, 11, 'lutff_5/lout')

wire n831;
// (7, 12, 'lutff_1/lout')

wire n832;
// (2, 8, 'lutff_5/lout')

wire n833;
// (5, 4, 'lutff_4/lout')

wire n834;
// (6, 8, 'lutff_6/lout')

wire n835;
// (4, 8, 'lutff_7/lout')

wire n836;
// (7, 4, 'lutff_6/lout')

wire n837;
// (7, 13, 'lutff_2/lout')

wire n838;
// (5, 5, 'lutff_5/lout')

wire n839;
// (9, 5, 'lutff_0/lout')

wire n840;
// (2, 12, 'lutff_2/lout')

wire n841;
// (7, 5, 'lutff_7/lout')

wire n842;
// (4, 12, 'lutff_4/lout')

wire n843;
// (6, 7, 'lutff_1/lout')

wire n844;
// (8, 7, 'lutff_3/lout')

wire n845;
// (5, 8, 'lutff_6/lout')

wire n846;
// (9, 8, 'lutff_1/lout')

wire n847;
// (4, 15, 'lutff_5/lout')

wire n848;
// (7, 11, 'lutff_4/lout')

wire n849;
// (4, 7, 'lutff_1/lout')

wire n850;
// (8, 11, 'lutff_0/lout')

wire n851;
// (6, 11, 'lutff_7/lout')

wire n852;
// (11, 6, 'lutff_7/lout')

wire n853;
// (11, 9, 'lutff_3/lout')

wire n854;
// (5, 12, 'lutff_3/lout')

wire n855;
// (7, 12, 'lutff_5/lout')

wire n856;
// (6, 8, 'lutff_1/lout')

wire n857;
// (4, 8, 'lutff_2/lout')

wire n858;
// (7, 4, 'lutff_1/lout')

wire n859;
// (8, 8, 'lutff_3/lout')

wire n860;
// (11, 10, 'lutff_4/lout')

wire n861;
// (5, 5, 'lutff_0/lout')

wire n862;
// (7, 5, 'lutff_2/lout')

wire n863;
// (9, 5, 'lutff_4/lout')

wire n864;
// (2, 4, 'lutff_2/lout')

wire n865;
// (4, 11, 'lutff_3/lout')

wire n866;
// (6, 15, 'lutff_0/lout')

wire n867;
// (6, 7, 'lutff_5/lout')

wire n868;
// (8, 7, 'lutff_7/lout')

wire n869;
// (11, 13, 'lutff_5/lout')

wire n870;
// (5, 8, 'lutff_1/lout')

wire n871;
// (4, 15, 'lutff_0/lout')

wire n872;
// (9, 8, 'lutff_5/lout')

wire n873;
// (5, 11, 'lutff_6/lout')

wire n874;
// (2, 7, 'lutff_3/lout')

wire n875;
// (4, 7, 'lutff_5/lout')

wire n876;
// (6, 11, 'lutff_2/lout')

wire n877;
// (8, 11, 'lutff_4/lout')

wire n878;
// (11, 9, 'lutff_7/lout')

wire n879;
// (7, 12, 'lutff_0/lout')

wire n880;
// (5, 4, 'lutff_3/lout')

wire n881;
// (4, 8, 'lutff_6/lout')

wire n882;
// (7, 4, 'lutff_5/lout')

wire n883;
// (6, 3, 'lutff_3/lout')

wire n884;
// (8, 14, 'lutff_5/lout')

wire n885;
// (7, 15, 'lutff_1/lout')

wire n886;
// (5, 7, 'lutff_4/lout')

wire n887;
// (6, 15, 'lutff_4/lout')

wire n888;
// (7, 7, 'lutff_6/lout')

wire n889;
// (4, 3, 'lutff_3/lout')

wire n890;
// (6, 7, 'lutff_0/lout')

wire n891;
// (4, 14, 'lutff_3/lout')

wire n892;
// (8, 7, 'lutff_2/lout')

wire n893;
// (11, 13, 'lutff_0/out')

wire n894;
// (11, 13, 'lutff_0/lout')

wire n895;
// (11, 13, 'carry_in_mux')

// Carry-In for (11 13)
assign n895 = 1;

wire n896;
// (11, 5, 'lutff_5/lout')

wire n897;
// (5, 8, 'lutff_5/lout')

wire n898;
// (9, 8, 'lutff_0/lout')

wire n899;
// (2, 15, 'lutff_2/lout')

wire n900;
// (5, 11, 'lutff_1/lout')

wire n901;
// (4, 15, 'lutff_4/lout')

wire n902;
// (7, 11, 'lutff_3/lout')

wire n903;
// (4, 7, 'lutff_0/lout')

wire n904;
// (2, 7, 'lutff_7/lout')

wire n905;
// (11, 6, 'lutff_6/lout')

wire n906;
// (11, 9, 'lutff_2/lout')

wire n907;
// (7, 12, 'lutff_4/lout')

wire n908;
// (4, 8, 'lutff_1/lout')

wire n909;
// (7, 4, 'lutff_0/lout')

wire n910;
// (8, 14, 'lutff_0/lout')

wire n911;
// (8, 3, 'lutff_0/lout')

wire n912;
// (6, 3, 'lutff_7/lout')

wire n913;
// (6, 14, 'lutff_7/lout')

wire n914;
// (4, 11, 'lutff_2/lout')

wire n915;
// (7, 7, 'lutff_1/lout')

wire n916;
// (9, 4, 'lutff_7/lout')

wire n917;
// (9, 7, 'lutff_3/lout')

wire n918;
// (4, 3, 'lutff_7/lout')

wire n919;
// (6, 7, 'lutff_4/lout')

wire n920;
// (8, 7, 'lutff_6/lout')

wire n921;
// (11, 13, 'lutff_4/lout')

wire n922;
// (11, 5, 'lutff_0/lout')

wire n923;
// (5, 8, 'lutff_0/lout')

wire n924;
// (9, 8, 'lutff_4/lout')

wire n925;
// (2, 15, 'lutff_6/lout')

wire n926;
// (2, 7, 'lutff_2/lout')

wire n927;
// (11, 6, 'lutff_1/lout')

wire n928;
// (5, 14, 'lutff_7/lout')

wire n929;
// (6, 10, 'lutff_5/lout')

wire n930;
// (11, 9, 'lutff_6/lout')

wire n931;
// (8, 10, 'lutff_7/lout')

wire n932;
// (9, 11, 'lutff_5/lout')

wire n933;
// (5, 3, 'lutff_6/lout')

wire n934;
// (4, 10, 'lutff_5/lout')

wire n935;
// (6, 14, 'lutff_2/lout')

wire n936;
// (6, 3, 'lutff_2/lout')

wire n937;
// (8, 14, 'lutff_4/lout')

wire n938;
// (8, 3, 'lutff_4/lout')

wire n939;
// (7, 15, 'lutff_0/lout')

wire n940;
// (11, 4, 'lutff_3/lout')

wire n941;
// (5, 15, 'lutff_7/lout')

wire n942;
// (5, 7, 'lutff_3/lout')

wire n943;
// (4, 11, 'lutff_6/lout')

wire n944;
// (7, 7, 'lutff_5/lout')

wire n945;
// (4, 3, 'lutff_2/lout')

wire n946;
// (4, 14, 'lutff_2/lout')

wire n947;
// (9, 7, 'lutff_7/lout')

wire n948;
// (8, 7, 'lutff_1/lout')

wire n949;
// (8, 6, 'lutff_5/lout')

wire n950;
// (5, 11, 'lutff_0/lout')

wire n951;
// (7, 11, 'lutff_2/lout')

wire n952;
// (7, 14, 'lutff_4/lout')

wire n953;
// (6, 10, 'lutff_0/lout')

wire n954;
// (11, 9, 'lutff_1/lout')

wire n955;
// (8, 10, 'lutff_2/lout')

wire n956;
// (6, 13, 'lutff_5/lout')

wire n957;
// (9, 11, 'lutff_0/lout')

wire n958;
// (5, 3, 'lutff_1/lout')

wire n959;
// (7, 3, 'lutff_3/lout')

wire n960;
// (9, 3, 'lutff_5/lout')

wire n961;
// (5, 6, 'lutff_6/lout')

wire n962;
// (6, 14, 'lutff_6/lout')

wire n963;
// (6, 6, 'lutff_2/lout')

wire n964;
// (5, 15, 'lutff_2/lout')

wire n965;
// (7, 15, 'lutff_4/lout')

wire n966;
// (7, 7, 'lutff_0/lout')

wire n967;
// (9, 4, 'lutff_6/lout')

wire n968;
// (5, 7, 'lutff_7/lout')

wire n969;
// (9, 7, 'lutff_2/lout')

wire n970;
// (11, 13, 'lutff_3/lout')

wire n971;
// (6, 9, 'lutff_3/lout')

wire n972;
// (8, 9, 'lutff_5/lout')

wire n973;
// (9, 14, 'lutff_1/lout')

wire n974;
// (4, 6, 'lutff_7/lout')

wire n975;
// (6, 10, 'lutff_4/lout')

wire n976;
// (6, 13, 'lutff_0/lout')

wire n977;
// (8, 10, 'lutff_6/lout')

wire n978;
// (9, 11, 'lutff_4/lout')

wire n979;
// (5, 3, 'lutff_5/lout')

wire n980;
// (5, 6, 'lutff_1/lout')

wire n981;
// (8, 14, 'lutff_3/lout')

wire n982;
// (8, 13, 'lutff_7/lout')

wire n983;
// (9, 4, 'lutff_1/lout')

wire n984;
// (5, 7, 'lutff_2/lout')

wire n985;
// (7, 7, 'lutff_4/lout')

wire n986;
// (4, 3, 'lutff_1/lout')

wire n987;
// (4, 14, 'lutff_1/out')

wire n988;
// (4, 14, 'lutff_1/lout')

wire n989;
// (9, 7, 'lutff_6/lout')

wire n990;
// (5, 10, 'lutff_4/lout')

wire n991;
// (7, 10, 'lutff_6/lout')

wire n992;
// (8, 6, 'lutff_4/lout')

wire n993;
// (8, 9, 'lutff_0/lout')

wire n994;
// (6, 9, 'lutff_7/lout')

wire n995;
// (7, 14, 'lutff_3/lout')

wire n996;
// (8, 10, 'lutff_1/lout')

wire n997;
// (6, 13, 'lutff_4/lout')

wire n998;
// (7, 3, 'lutff_2/lout')

wire n999;
// (9, 3, 'lutff_4/lout')

wire n1000;
// (2, 10, 'lutff_6/lout')

wire n1001;
// (5, 6, 'lutff_5/lout')

wire n1002;
// (7, 6, 'lutff_4/lout')

wire n1003;
// (11, 12, 'lutff_1/lout')

wire n1004;
// (8, 13, 'lutff_2/lout')

wire n1005;
// (5, 9, 'lutff_7/lout')

wire n1006;
// (1, 12, 'lutff_0/lout')

wire n1007;
// (6, 5, 'lutff_5/lout')

wire n1008;
// (8, 5, 'lutff_7/lout')

wire n1009;
// (7, 10, 'lutff_1/lout')

wire n1010;
// (9, 10, 'lutff_3/lout')

wire n1011;
// (6, 9, 'lutff_2/lout')

wire n1012;
// (8, 9, 'lutff_4/lout')

wire n1013;
// (11, 7, 'lutff_7/lout')

wire n1014;
// (2, 6, 'lutff_4/lout')

wire n1015;
// (12, 7, 'lutff_3/lout')

wire n1016;
// (7, 14, 'lutff_7/lout')

wire n1017;
// (6, 12, 'lutff_3/lout')

wire n1018;
// (8, 12, 'lutff_5/lout')

wire n1019;
// (5, 6, 'lutff_0/lout')

wire n1020;
// (9, 6, 'lutff_1/lout')

wire n1021;
// (5, 9, 'lutff_2/lout')

wire n1022;
// (7, 9, 'lutff_4/lout')

wire n1023;
// (6, 5, 'lutff_0/lout')

wire n1024;
// (8, 13, 'lutff_6/lout')

wire n1025;
// (11, 11, 'lutff_0/lout')

wire n1026;
// (9, 9, 'lutff_6/lout')

wire n1027;
// (8, 5, 'lutff_2/lout')

wire n1028;
// (7, 10, 'lutff_5/lout')

wire n1029;
// (9, 10, 'lutff_7/lout')

wire n1030;
// (6, 9, 'lutff_6/lout')

wire n1031;
// (4, 9, 'lutff_7/lout')

wire n1032;
// (11, 7, 'lutff_2/lout')

wire n1033;
// (4, 6, 'lutff_1/lout')

wire n1034;
// (7, 14, 'lutff_2/lout')

wire n1035;
// (7, 13, 'lutff_6/lout')

wire n1036;
// (11, 8, 'lutff_3/lout')

wire n1037;
// (8, 12, 'lutff_0/lout')

wire n1038;
// (2, 12, 'lutff_6/lout')

wire n1039;
// (6, 12, 'lutff_7/lout')

wire n1040;
// (6, 4, 'lutff_3/lout')

wire n1041;
// (8, 4, 'lutff_5/lout')

wire n1042;
// (7, 6, 'lutff_3/lout')

wire n1043;
// (9, 6, 'lutff_5/lout')

wire n1044;
// (2, 13, 'lutff_7/lout')

wire n1045;
// (5, 9, 'lutff_6/lout')

wire n1046;
// (8, 13, 'lutff_1/lout')

wire n1047;
// (9, 9, 'lutff_1/lout')

wire n1048;
// (6, 5, 'lutff_4/lout')

wire n1049;
// (8, 5, 'lutff_6/lout')

wire n1050;
// (11, 11, 'lutff_4/lout')

wire n1051;
// (9, 10, 'lutff_2/lout')

wire n1052;
// (8, 9, 'lutff_3/lout')

wire n1053;
// (11, 7, 'lutff_6/lout')

wire n1054;
// (8, 8, 'lutff_7/lout')

wire n1055;
// (7, 13, 'lutff_1/lout')

wire n1056;
// (9, 13, 'lutff_3/lout')

wire n1057;
// (2, 12, 'lutff_1/lout')

wire n1058;
// (7, 5, 'lutff_6/lout')

wire n1059;
// (6, 12, 'lutff_2/lout')

wire n1060;
// (4, 12, 'lutff_3/lout')

wire n1061;
// (8, 12, 'lutff_4/lout')

wire n1062;
// (8, 4, 'lutff_0/lout')

wire n1063;
// (6, 4, 'lutff_7/lout')

wire n1064;
// (9, 6, 'lutff_0/lout')

wire n1065;
// (5, 9, 'lutff_1/lout')

wire n1066;
// (7, 6, 'lutff_7/lout')

wire n1067;
// (7, 9, 'lutff_3/lout')

wire n1068;
// (8, 13, 'lutff_5/lout')

wire n1069;
// (9, 9, 'lutff_5/lout')

wire n1070;
// (8, 5, 'lutff_1/lout')

wire n1071;
// (6, 11, 'lutff_6/lout')

wire n1072;
// (6, 8, 'lutff_0/lout')

wire n1073;
// (8, 8, 'lutff_2/lout')

wire n1074;
// (5, 4, 'lutff_7/lout')

wire n1075;
// (7, 13, 'lutff_5/lout')

wire n1076;
// (7, 5, 'lutff_1/lout')

wire n1077;
// (12, 9, 'lutff_6/lout')

wire n1078;
// (9, 5, 'lutff_3/lout')

wire n1079;
// (6, 12, 'lutff_6/lout')

wire n1080;
// (4, 12, 'lutff_7/lout')

wire n1081;
// (6, 4, 'lutff_2/lout')

wire n1082;
// (8, 4, 'lutff_4/lout')

wire n1083;
// (7, 6, 'lutff_2/lout')

wire n1084;
// (9, 6, 'lutff_4/lout')

wire n1085;
// (5, 9, 'lutff_5/lout')

wire n1086;
// (9, 9, 'lutff_0/lout')

wire n1087;
// (2, 5, 'lutff_2/lout')

wire n1088;
// (7, 9, 'lutff_7/lout')

wire n1089;
// (6, 11, 'lutff_1/lout')

wire n1090;
// (8, 11, 'lutff_3/lout')

assign n663  = /* LUT    4 14  0 */ 1'b0;
assign n693  = /* LUT   11 13  1 */ 1'b0;
assign n894  = /* LUT   11 13  0 */ 1'b0;
assign n988  = /* LUT    4 14  1 */ 1'b0;
assign n547  = /* LUT    5 12  6 */ n184;
assign n548  = /* LUT    9 12  1 */ (n371 ? (n188 ? (n455 ? 1'b0 : !n433) : 1'b0) : 1'b0);
assign n549  = /* LUT    5  4  2 */ (n139 ? (n160 ? (n84 ? 1'b1 : n189) : (n84 ? n189 : 1'b1)) : (n160 ? (n84 ? 1'b0 : !n189) : (n84 ? !n189 : 1'b0)));
assign n550  = /* LUT    4  8  5 */ n108;
assign n551  = /* LUT    8  8  6 */ (n23 ? (n409 ? (n321 ? 1'b1 : n189) : (n321 ? n189 : 1'b1)) : (n409 ? (n321 ? 1'b0 : !n189) : (n321 ? !n189 : 1'b0)));
assign n552  = /* LUT    7  4  4 */ n304;
assign n553  = /* LUT    7 13  0 */ (n365 ? (n276 ? !n280 : n280) : 1'b0);
assign n554  = /* LUT    9 13  2 */ (n512 ? (n455 ? !n371 : n371) : 1'b0);
assign n555  = /* LUT    5  5  3 */ n152;
assign n556  = /* LUT    6 12  1 */ (n268 ? 1'b0 : !n265);
assign n557  = /* LUT    7  5  5 */ n312;
assign n558  = /* LUT    4 12  2 */ (n119 ? (n38 ? 1'b1 : (n58 ? 1'b1 : n52)) : 1'b0);
assign n559  = /* LUT    8 12  3 */ (n356 ? (n364 ? (n2 ? !n435 : 1'b0) : (n2 ? n435 : 1'b1)) : (n364 ? (n2 ? n435 : 1'b1) : (n2 ? !n435 : 1'b0)));
assign n560  = /* LUT    6 15  3 */ (n281 ? n288 : !n288);
assign n561  = /* LUT    5  9  0 */ (n106 ? n53 : !n53);
assign n562  = /* LUT    9  9  4 */ (n499 ? (n478 ? !n416 : n416) : (n478 ? n416 : !n416));
assign n563  = /* LUT    5  8  4 */ n170;
assign n564  = /* LUT    7  8  6 */ (n10 ? (n15 ? !n20 : 1'b1) : (n15 ? n20 : 1'b0));
assign n565  = /* LUT    4 15  3 */ (n128 ? (n64 ? 1'b0 : (n39 ? 1'b1 : !n123)) : 1'b0);
assign n566  = /* LUT   11  6  5 */ n69;
assign n567  = /* LUT    8 11  7 */ (n352 ? (n201 ? 1'b0 : n353) : (n201 ? 1'b1 : n336));
assign n568  = /* LUT    5 12  1 */ (n91 ? (n38 ? 1'b0 : (n58 ? 1'b0 : !n52)) : 1'b0);
assign n569  = /* LUT    7 12  3 */ (n35 ? (n436 ? (n354 ? n195 : !n195) : (n354 ? !n195 : n195)) : 1'b0);
assign n570  = /* LUT    4  8  0 */ n97;
assign n571  = /* LUT    8  8  1 */ n413;
assign n572  = /* LUT    5  4  6 */ n153;
assign n573  = /* LUT    7 13  4 */ (n277 ? (n365 ? n122 : 1'b1) : (n365 ? (n122 ? n449 : !n449) : !n449));
assign n574  = /* LUT    7  5  0 */ (n68 ? (n7 ? 1'b1 : !n225) : (n7 ? 1'b0 : n229));
assign n575  = /* LUT    5  5  7 */ n147;
assign n576  = /* LUT    9  5  2 */ n476;
assign n577  = /* LUT    2 12  4 */ n27;
assign n578  = /* LUT    2  4  0 */ n66;
assign n579  = /* LUT    4 12  6 */ n90;
assign n580  = /* LUT    6 15  7 */ (n284 ? (n274 ? (n285 ? 1'b0 : n286) : (n285 ? n286 : 1'b0)) : (n274 ? (n285 ? 1'b1 : !n286) : (n285 ? !n286 : 1'b1)));
assign n581  = /* LUT    6  7  3 */ (n7 ? (n107 ? n240 : n102) : n240);
assign n582  = /* LUT    7  8  1 */ n327;
assign n583  = /* LUT    5 11  4 */ (n185 ? (n38 ? 1'b0 : (n58 ? 1'b0 : !n52)) : 1'b0);
assign n584  = /* LUT    4 15  7 */ (n52 ? (n131 ? 1'b0 : (n123 ? !n39 : 1'b1)) : (n123 ? !n39 : 1'b1));
assign n585  = /* LUT    7 11  6 */ (n353 ? (n352 ? (n336 ? !n201 : 1'b0) : (n336 ? n201 : !n201)) : (n352 ? (n336 ? n201 : 1'b1) : n201));
assign n586  = /* LUT    4  7  3 */ n93;
assign n587  = /* LUT   11  6  0 */ (n107 ? (n7 ? 1'b1 : !n485) : (n7 ? !n484 : 1'b1));
assign n588  = /* LUT    8 11  2 */ (n275 ? (n429 ? 1'b1 : n344) : (n429 ? (n347 ? n344 : !n344) : n347));
assign n589  = /* LUT   11  9  5 */ (n406 ? (n15 ? !n527 : 1'b1) : (n15 ? n527 : 1'b0));
assign n590  = /* LUT    5 12  5 */ (n56 ? (n204 ? (n195 ? !n35 : 1'b1) : (n195 ? 1'b1 : !n35)) : (n204 ? (n195 ? n35 : 1'b0) : (n195 ? 1'b0 : n35)));
assign n591  = /* LUT    7 12  7 */ (n2 ? (n437 ? (n188 ? !n433 : 1'b0) : 1'b0) : 1'b0);
assign n592  = /* LUT    5  4  1 */ n141;
assign n593  = /* LUT    6  8  3 */ (n42 ? n245 : n246);
assign n594  = /* LUT    4  8  4 */ (n106 ? n33 : !n33);
assign n595  = /* LUT    7  4  3 */ n295;
assign n596  = /* LUT    8  8  5 */ n410;
assign n597  = /* LUT    6  3  1 */ (n42 ? n213 : n212);
assign n598  = /* LUT    6 14  1 */ (n273 ? n278 : !n278);
assign n599  = /* LUT    8  3  3 */ (n101 ? n460 : !n65);
assign n600  = /* LUT    6  6  6 */ n231;
assign n601  = /* LUT    4 11  5 */ n194;
assign n602  = /* LUT    6 15  2 */ (n288 ? (n289 ? (n287 ? !n132 : 1'b0) : (n287 ? 1'b0 : !n132)) : (n289 ? (n287 ? 1'b0 : !n132) : (n287 ? !n132 : 1'b0)));
assign n603  = /* LUT    8  7  0 */ (n169 ? (n42 ? n405 : n486) : (n42 ? !n405 : !n486));
assign n604  = /* LUT    6  7  7 */ n238;
assign n605  = /* LUT   11 13  7 */ (n544 ? !n371 : n371);
assign n606  = /* LUT    5  8  3 */ n172;
assign n607  = /* LUT    7  8  5 */ n330;
assign n608  = /* LUT    4 15  2 */ (n127 ? (n126 ? 1'b0 : (n125 ? 1'b0 : !n124)) : 1'b0);
assign n609  = /* LUT    9  8  7 */ n491;
assign n610  = /* LUT    7 11  1 */ (n201 ? (n353 ? 1'b0 : (n352 ? 1'b1 : n336)) : (n353 ? n336 : (n352 ? n336 : 1'b1)));
assign n611  = /* LUT    4  7  7 */ n86;
assign n612  = /* LUT    6 11  4 */ (n30 ? 1'b0 : !n266);
assign n613  = /* LUT    8 11  6 */ (n201 ? (n353 ? (n336 ? n352 : 1'b1) : (n336 ? 1'b1 : n352)) : (n353 ? n352 : 1'b0));
assign n614  = /* LUT   11  6  4 */ n516;
assign n615  = /* LUT   11  9  0 */ (n257 ? (n42 ? n525 : n524) : (n42 ? !n525 : !n524));
assign n616  = /* LUT    5 12  0 */ (n200 ? (n38 ? 1'b1 : (n58 ? 1'b1 : n52)) : 1'b0);
assign n617  = /* LUT    7 12  2 */ (n35 ? (n349 ? (n354 ? n195 : !n195) : (n354 ? !n195 : n195)) : 1'b0);
assign n618  = /* LUT    5  4  5 */ n9;
assign n619  = /* LUT    2 11  2 */ (n60 ? (n38 ? 1'b1 : (n58 ? 1'b1 : n52)) : 1'b0);
assign n620  = /* LUT    7  4  7 */ n301;
assign n621  = /* LUT    6  3  5 */ (n10 ? (n8 ? (n214 ? n15 : 1'b0) : (n214 ? !n15 : 1'b1)) : (n8 ? (n214 ? !n15 : 1'b1) : (n214 ? n15 : 1'b0)));
assign n622  = /* LUT    6 14  5 */ (n274 ? (n36 ? !n357 : 1'b1) : (n282 ? (n36 ? !n357 : 1'b1) : (n36 ? n357 : 1'b0)));
assign n623  = /* LUT    8 14  7 */ (n36 ? (n77 ? 1'b0 : !n451) : (n77 ? (n452 ? !n451 : n451) : !n452));
assign n624  = /* LUT    6  6  1 */ (n90 ? (n42 ? n243 : n250) : (n42 ? !n243 : !n250));
assign n625  = /* LUT    8  3  7 */ n381;
assign n626  = /* LUT    4 11  0 */ (n114 ? !n28 : !n109);
assign n627  = /* LUT    5  7  6 */ n18;
assign n628  = /* LUT    9  7  1 */ (n107 ? (n7 ? !n248 : 1'b1) : (n7 ? !n482 : 1'b0));
assign n629  = /* LUT    2  3  3 */ n43;
assign n630  = /* LUT    4 14  5 */ (n127 ? 1'b0 : (n35 ? (n123 ? 1'b1 : n205) : 1'b1));
assign n631  = /* LUT    6  7  2 */ (n107 ? (n7 ? n161 : n102) : n161);
assign n632  = /* LUT   11 13  2 */ (n539 ? !n530 : n530);
assign n633  = /* LUT    5  8  7 */ (n106 ? (n167 ? (n15 ? !n162 : 1'b1) : (n15 ? n162 : 1'b0)) : (n167 ? (n15 ? n162 : 1'b0) : (n15 ? !n162 : 1'b1)));
assign n634  = /* LUT    9  8  2 */ n490;
assign n635  = /* LUT    5 11  3 */ (n111 ? (n38 ? 1'b1 : (n58 ? 1'b1 : n52)) : 1'b0);
assign n636  = /* LUT    2  7  0 */ (n42 ? n70 : n49);
assign n637  = /* LUT    4 15  6 */ (n127 ? (n126 ? (n125 ? 1'b0 : !n124) : 1'b0) : 1'b0);
assign n638  = /* LUT    4  7  2 */ n92;
assign n639  = /* LUT    8 11  1 */ (n275 ? (n429 ? 1'b1 : n347) : (n429 ? n344 : (n347 ? n344 : !n344)));
assign n640  = /* LUT    6 10  3 */ n260;
assign n641  = /* LUT   11  9  4 */ (n406 ? (n15 ? !n526 : 1'b1) : (n15 ? n526 : 1'b0));
assign n642  = /* LUT    8 10  5 */ (n422 ? (n432 ? (n415 ? 1'b1 : !n345) : (n415 ? 1'b0 : n345)) : (n415 ? 1'b0 : n345));
assign n643  = /* LUT    5  4  0 */ (n145 ? (n146 ? (n83 ? 1'b1 : n189) : (n83 ? n189 : 1'b1)) : (n146 ? (n83 ? 1'b0 : !n189) : (n83 ? !n189 : 1'b0)));
assign n644  = /* LUT    7  4  2 */ n303;
assign n645  = /* LUT    9 11  3 */ (n421 ? (n416 ? n348 : !n348) : 1'b0);
assign n646  = /* LUT    7  3  6 */ n298;
assign n647  = /* LUT    4 10  3 */ n169;
assign n648  = /* LUT    6  3  0 */ (n184 ? (n42 ? n216 : n211) : (n42 ? !n216 : !n211));
assign n649  = /* LUT    6 14  0 */ (n278 ? (n133 ? !n273 : 1'b0) : (n133 ? (n273 ? !n77 : n77) : n77));
assign n650  = /* LUT    8 14  2 */ (n362 ? (n363 ? (n132 ? n208 : !n208) : n132) : (n363 ? n208 : (n132 ? n208 : !n208)));
assign n651  = /* LUT    8  3  2 */ n383;
assign n652  = /* LUT    6  6  5 */ n221;
assign n653  = /* LUT   11 12  5 */ (rst ? 1'b1 : (n203 ? 1'b1 : n39));
assign n654  = /* LUT    9  4  0 */ (n463 ? (n313 ? (n444 ? 1'b1 : n189) : (n444 ? n189 : 1'b1)) : (n313 ? (n444 ? 1'b0 : !n189) : (n444 ? !n189 : 1'b0)));
assign n655  = /* LUT    5  7  1 */ n236;
assign n656  = /* LUT    7 15  7 */ (n373 ? 1'b0 : (n374 ? 1'b0 : (n363 ? n290 : 1'b1)));
assign n657  = /* LUT    4 11  4 */ n115;
assign n658  = /* LUT    6 15  1 */ (n288 ? (n289 ? !n287 : n287) : (n289 ? n287 : !n287));
assign n659  = /* LUT    7  7  3 */ n324;
assign n660  = /* LUT    4  3  0 */ n81;
assign n661  = /* LUT    9  7  5 */ (n7 ? (n107 ? n482 : n248) : n482);
assign n665  = /* LUT   11 13  6 */ (n543 ? !n455 : n455);
assign n666  = /* LUT   12 12  0 */ !rst;
assign n667  = /* LUT    5  8  2 */ n175;
assign n668  = /* LUT    4 15  1 */ (n127 ? (n126 ? (n125 ? n124 : 1'b0) : 1'b0) : 1'b0);
assign n669  = /* LUT    4  4  1 */ (n146 ? !n83 : n83);
assign n670  = /* LUT    7 11  0 */ (n352 ? (n336 ? n353 : (n353 ? 1'b0 : n201)) : (n336 ? n353 : (n353 ? 1'b1 : !n201)));
assign n671  = /* LUT    4  7  6 */ n169;
assign n672  = /* LUT   11  6  3 */ n517;
assign n673  = /* LUT    8 10  0 */ (n334 ? (n432 ? n415 : 1'b1) : (n432 ? (n415 ? !n431 : n431) : n431));
assign n674  = /* LUT    6 10  7 */ n262;
assign n675  = /* LUT    6 13  3 */ (n113 ? (n75 ? !n74 : n74) : (n75 ? n74 : !n74));
assign n676  = /* LUT    7  3  1 */ n294;
assign n677  = /* LUT    9 11  7 */ (n426 ? (n504 ? n509 : !n509) : (n504 ? !n509 : n509));
assign n678  = /* LUT    9  3  3 */ n459;
assign n679  = /* LUT    5  6  4 */ (n166 ? (n15 ? !n154 : 1'b1) : (n15 ? n154 : 1'b0));
assign n680  = /* LUT    6  3  4 */ (n8 ? (n15 ? !n216 : 1'b1) : (n15 ? n216 : 1'b0));
assign n681  = /* LUT    6 14  4 */ (n282 ? n133 : !n133);
assign n682  = /* LUT    8  3  6 */ (n7 ? (n107 ? n376 : n460) : n376);
assign n683  = /* LUT    8 14  6 */ (n357 ? (n278 ? n452 : 1'b1) : (n278 ? (n452 ? n451 : !n451) : n451));
assign n684  = /* LUT    5 15  0 */ (n205 ? (n129 ? !rst : 1'b0) : 1'b0);
assign n685  = /* LUT    7 15  2 */ (n274 ? n285 : !n285);
assign n686  = /* LUT    9  4  4 */ n465;
assign n687  = /* LUT    5  7  5 */ n89;
assign n688  = /* LUT    9  7  0 */ (n397 ? (n159 ? (n493 ? !n472 : 1'b1) : (n493 ? n472 : 1'b0)) : (n159 ? (n493 ? n472 : 1'b0) : (n493 ? !n472 : 1'b1)));
assign n689  = /* LUT    7  7  7 */ (n7 ? (n107 ? n328 : n314) : n328);
assign n690  = /* LUT    4  3  4 */ n137;
assign n691  = /* LUT    4 14  4 */ (n127 ? (n126 ? 1'b0 : !n130) : (n126 ? !n130 : 1'b0));
assign n694  = /* LUT   11  5  6 */ n515;
assign n695  = /* LUT    6  9  1 */ (n42 ? n251 : n249);
assign n696  = /* LUT    8  6  7 */ n398;
assign n697  = /* LUT    7 14  6 */ (n362 ? (n132 ? (n363 ? 1'b0 : n208) : n363) : (n132 ? (n363 ? 1'b0 : !n208) : 1'b1));
assign n698  = /* LUT    8 10  4 */ (n432 ? (n498 ? (n416 ? !n345 : 1'b1) : (n416 ? n345 : 1'b0)) : (n416 ? !n345 : 1'b1));
assign n699  = /* LUT    6 13  7 */ (n113 ? (n74 ? !n198 : n198) : (n74 ? n198 : !n198));
assign n700  = /* LUT    6  2  7 */ n214;
assign n701  = /* LUT    9 11  2 */ (n159 ? (n497 ? !n506 : 1'b0) : (n497 ? 1'b0 : !n506));
assign n702  = /* LUT    5  3  3 */ n138;
assign n703  = /* LUT    4 10  2 */ n108;
assign n704  = /* LUT    8  3  1 */ (n107 ? (n7 ? !n460 : 1'b1) : (n7 ? !n376 : 1'b0));
assign n705  = /* LUT    8 14  1 */ (n362 ? (n363 ? (n132 ? n208 : !n208) : (n132 ? 1'b0 : n208)) : (n363 ? (n132 ? !n208 : 1'b0) : 1'b1));
assign n706  = /* LUT    6  6  4 */ n244;
assign n707  = /* LUT   11 12  4 */ (n534 ? 1'b0 : (n76 ? 1'b0 : (n530 ? 1'b0 : !n34)));
assign n708  = /* LUT    5  7  0 */ (n108 ? (n42 ? n162 : n46) : (n42 ? !n162 : !n46));
assign n709  = /* LUT    7 15  6 */ (n291 ? (n292 ? (n453 ? 1'b0 : !n132) : 1'b0) : (n292 ? 1'b0 : (n453 ? !n132 : 1'b0)));
assign n710  = /* LUT    7  7  2 */ n326;
assign n711  = /* LUT    9  7  4 */ n494;
assign n712  = /* LUT    5 10  2 */ n91;
assign n713  = /* LUT    7 10  4 */ (n423 ? (n346 ? (n264 ? n342 : !n342) : n342) : (n346 ? n264 : 1'b0));
assign n714  = /* LUT    8  6  2 */ (n396 ? (n7 ? 1'b1 : !n384) : (n7 ? 1'b0 : n47));
assign n715  = /* LUT    9 10  6 */ (n264 ? (n423 ? 1'b0 : !n503) : (n423 ? !n503 : 1'b0));
assign n716  = /* LUT    6  9  5 */ (n8 ? (n242 ? (n24 ? !n15 : 1'b1) : (n24 ? n15 : 1'b0)) : (n242 ? (n24 ? n15 : 1'b0) : (n24 ? !n15 : 1'b1)));
assign n717  = /* LUT    8  9  7 */ (n428 ? (n419 ? (n337 ? n417 : !n417) : (n337 ? !n417 : n417)) : (n419 ? (n337 ? !n417 : n417) : (n337 ? n417 : !n417)));
assign n718  = /* LUT    7 14  1 */ (n362 ? (n208 ? 1'b0 : !n132) : (n208 ? 1'b1 : n363));
assign n719  = /* LUT   12  7  6 */ n535;
assign n720  = /* LUT    6 10  6 */ n258;
assign n721  = /* LUT    6 13  2 */ (n74 ? !n198 : n198);
assign n722  = /* LUT    9 11  6 */ (n505 ? (n159 ? (n497 ? 1'b0 : n506) : (n497 ? n506 : 1'b0)) : (n159 ? (n497 ? 1'b1 : !n506) : (n497 ? !n506 : 1'b1)));
assign n723  = /* LUT    7  3  0 */ n305;
assign n724  = /* LUT    5  3  7 */ n136;
assign n725  = /* LUT    5  6  3 */ (n42 ? n156 : n13);
assign n726  = /* LUT    4 10  6 */ n176;
assign n727  = /* LUT    8 13  0 */ (n450 ? (n355 ? (n446 ? n441 : !n441) : (n446 ? !n441 : n441)) : (n355 ? (n446 ? !n441 : n441) : (n446 ? n441 : !n441)));
assign n728  = /* LUT    6  5  3 */ (n107 ? (n7 ? n225 : n226) : n225);
assign n729  = /* LUT    8  5  5 */ (n107 ? (n7 ? n384 : n392) : n384);
assign n730  = /* LUT    5 10  6 */ (n173 ? (n33 ? n189 : 1'b1) : (n33 ? !n189 : 1'b0));
assign n731  = /* LUT    9 10  1 */ (n159 ? (n478 ? (n264 ? n334 : !n334) : (n264 ? !n334 : n334)) : (n478 ? (n264 ? !n334 : n334) : (n264 ? n334 : !n334)));
assign n732  = /* LUT    6  9  0 */ (n42 ? n252 : n25);
assign n733  = /* LUT    8  6  6 */ (n241 ? (n88 ? n189 : 1'b1) : (n88 ? !n189 : 1'b0));
assign n734  = /* LUT   11  7  5 */ n519;
assign n735  = /* LUT   12  7  1 */ n73;
assign n736  = /* LUT    6 10  1 */ n261;
assign n737  = /* LUT    7 14  5 */ (n372 ? (n282 ? 1'b1 : n366) : (n282 ? 1'b0 : !n366));
assign n738  = /* LUT    8 10  3 */ (n496 ? !n334 : n334);
assign n739  = /* LUT    6 13  6 */ (n122 ? (n277 ? (n269 ? n276 : !n276) : n269) : (n277 ? 1'b0 : n276));
assign n740  = /* LUT    9 11  1 */ (n501 ? (n509 ? !n508 : n508) : (n509 ? n508 : !n508));
assign n741  = /* LUT    5  3  2 */ n135;
assign n742  = /* LUT    7  3  4 */ n296;
assign n743  = /* LUT    9  3  6 */ n457;
assign n744  = /* LUT    5  6  7 */ (n42 ? n157 : n155);
assign n745  = /* LUT    7  6  6 */ n230;
assign n746  = /* LUT   11 12  3 */ (rst ? 1'b1 : (n531 ? n533 : 1'b0));
assign n747  = /* LUT    8 13  4 */ (n35 ? (n513 ? n447 : !n447) : 1'b0);
assign n748  = /* LUT    8  5  0 */ n394;
assign n749  = /* LUT    6  5  7 */ n222;
assign n750  = /* LUT   11 11  7 */ (n76 ? (n34 ? 1'b1 : n534) : (n34 ? n534 : 1'b1));
assign n751  = /* LUT    5 10  1 */ n51;
assign n752  = /* LUT    7 10  3 */ (n348 ? (n346 ? n159 : 1'b1) : (n346 ? (n159 ? n342 : !n342) : !n342));
assign n753  = /* LUT    8  6  1 */ (n107 ? (n7 ? !n392 : 1'b1) : (n7 ? !n391 : 1'b0));
assign n754  = /* LUT    9 10  5 */ (n264 ? !n334 : n334);
assign n755  = /* LUT    6  9  4 */ (n8 ? (n15 ? !n252 : 1'b1) : (n15 ? n252 : 1'b0));
assign n756  = /* LUT    4  9  5 */ n24;
assign n757  = /* LUT    8  9  6 */ (n430 ? (n420 ? (n428 ? n338 : !n338) : (n428 ? !n338 : n338)) : (n420 ? (n428 ? !n338 : n338) : (n428 ? n338 : !n338)));
assign n758  = /* LUT   11  7  0 */ (n42 ? n72 : n521);
assign n759  = /* LUT    7 14  0 */ (n375 ? (n274 ? 1'b1 : n366) : (n274 ? 1'b0 : !n366));
assign n760  = /* LUT   11  8  1 */ n255;
assign n761  = /* LUT    6 12  5 */ (n271 ? (n267 ? !n199 : n199) : (n267 ? n199 : !n199));
assign n762  = /* LUT    8 12  7 */ (n356 ? (n364 ? (n2 ? n438 : 1'b1) : (n2 ? !n438 : 1'b0)) : (n364 ? (n2 ? !n438 : 1'b0) : (n2 ? n438 : 1'b1)));
assign n763  = /* LUT    7  6  1 */ n318;
assign n764  = /* LUT    9  6  3 */ (n7 ? (n107 ? n484 : n477) : n484);
assign n765  = /* LUT    5  9  4 */ (n53 ? (n15 ? !n182 : 1'b1) : (n15 ? n182 : 1'b0));
assign n766  = /* LUT    4 13  7 */ (n4 ? (n123 ? 1'b1 : rst) : 1'b1);
assign n767  = /* LUT    2  5  1 */ n67;
assign n768  = /* LUT    7  9  6 */ (n307 ? (n377 ? (n159 ? !n234 : n234) : (n159 ? n234 : !n234)) : (n377 ? (n159 ? n234 : !n234) : (n159 ? !n234 : n234)));
assign n769  = /* LUT    6  5  2 */ n227;
assign n770  = /* LUT    8  5  4 */ n390;
assign n771  = /* LUT    5 10  5 */ (n263 ? (n242 ? !n202 : n202) : (n242 ? n202 : !n202));
assign n772  = /* LUT    9 10  0 */ (n416 ? (n397 ? 1'b0 : !n497) : (n397 ? (n497 ? !n334 : n334) : n334));
assign n773  = /* LUT    7 10  7 */ (n340 ? (n424 ? (n427 ? !n418 : n418) : (n427 ? n418 : !n418)) : (n424 ? (n427 ? n418 : !n418) : (n427 ? !n418 : n418)));
assign n774  = /* LUT    8  9  1 */ (n307 ? (n377 ? !n159 : n159) : (n377 ? n159 : !n159));
assign n775  = /* LUT   11  7  4 */ (n101 ? n248 : !n492);
assign n776  = /* LUT    4  6  3 */ n88;
assign n777  = /* LUT    5  5  2 */ n90;
assign n778  = /* LUT    6 12  0 */ (n268 ? (n190 ? 1'b0 : !n197) : (n190 ? !n265 : (n197 ? !n265 : n265)));
assign n779  = /* LUT    7  5  4 */ n310;
assign n780  = /* LUT    4 12  1 */ (n44 ? (n38 ? 1'b0 : (n58 ? 1'b0 : !n52)) : 1'b0);
assign n781  = /* LUT    8 12  2 */ (n371 ? (n188 ? 1'b1 : (n433 ? 1'b1 : n455)) : (n188 ? (n433 ? n455 : 1'b1) : 1'b1));
assign n782  = /* LUT    9  5  6 */ n469;
assign n783  = /* LUT    8  4  7 */ n385;
assign n784  = /* LUT    7  6  5 */ n315;
assign n785  = /* LUT    8 13  3 */ (n2 ? (n455 ? 1'b0 : !n188) : 1'b0);
assign n786  = /* LUT    7  9  1 */ (n419 ? n338 : !n338);
assign n787  = /* LUT    9  6  7 */ n473;
assign n788  = /* LUT    6  5  6 */ n224;
assign n789  = /* LUT    5 10  0 */ n185;
assign n790  = /* LUT    7 10  2 */ (n159 ? (n346 ? !n348 : 1'b0) : (n346 ? (n348 ? n343 : !n343) : !n343));
assign n791  = /* LUT    9 10  4 */ (n496 ? (n478 ? (n264 ? !n334 : 1'b0) : (n264 ? 1'b0 : !n334)) : (n478 ? (n264 ? 1'b0 : n334) : (n264 ? n334 : 1'b0)));
assign n792  = /* LUT    8  8  0 */ (n106 ? !n407 : n407);
assign n793  = /* LUT    2  8  6 */ n21;
assign n794  = /* LUT    6  8  7 */ (n333 ? !n242 : n242);
assign n795  = /* LUT    7 13  3 */ (n276 ? (n365 ? n280 : 1'b1) : (n365 ? (n280 ? !n370 : n370) : n370));
assign n796  = /* LUT    9 13  5 */ (n76 ? !n34 : n34);
assign n797  = /* LUT    5  5  6 */ n149;
assign n798  = /* LUT    9  5  1 */ n475;
assign n799  = /* LUT    6 12  4 */ (n271 ? (n269 ? !n199 : n199) : (n269 ? n199 : !n199));
assign n800  = /* LUT    4 12  5 */ (n117 ? (n118 ? 1'b1 : n31) : (n118 ? n116 : (n31 ? n116 : !n116)));
assign n801  = /* LUT    6  4  0 */ n143;
assign n802  = /* LUT    8 12  6 */ (n455 ? (n371 ? 1'b1 : (n188 ? 1'b1 : n433)) : (n371 ? n188 : 1'b1));
assign n803  = /* LUT    8  4  2 */ n387;
assign n804  = /* LUT    7  6  0 */ n317;
assign n805  = /* LUT    9  6  2 */ n467;
assign n806  = /* LUT    5  9  3 */ (n106 ? (n15 ? n177 : 1'b0) : (n15 ? !n177 : 1'b1));
assign n807  = /* LUT    7  9  5 */ (n307 ? (n377 ? (n159 ? !n322 : n322) : (n159 ? n322 : !n322)) : (n377 ? (n159 ? n322 : !n322) : (n159 ? !n322 : n322)));
assign n808  = /* LUT    6  5  1 */ n308;
assign n809  = /* LUT    8  5  3 */ n389;
assign n810  = /* LUT    5 12  4 */ (n196 ? 1'b0 : !n193);
assign n811  = /* LUT    7  1  6 */ !n42;
assign n812  = /* LUT    6  8  2 */ (n106 ? (n15 ? n245 : 1'b0) : (n15 ? !n245 : 1'b1));
assign n813  = /* LUT    7 12  6 */ (n35 ? (n350 ? (n195 ? !n361 : n361) : (n195 ? n361 : !n361)) : 1'b0);
assign n814  = /* LUT    4  8  3 */ n99;
assign n815  = /* LUT    8  8  4 */ (n409 ? (n406 ? n321 : !n321) : (n406 ? !n321 : n321));
assign n816  = /* LUT    2 11  6 */ n59;
assign n817  = /* LUT    9 13  0 */ (n2 ? (n433 ? !n188 : 1'b0) : 1'b0);
assign n818  = /* LUT    5  5  1 */ n150;
assign n819  = /* LUT    7 13  7 */ (n367 ? (n359 ? (n293 ? n441 : !n441) : (n293 ? !n441 : n441)) : (n359 ? (n293 ? !n441 : n441) : (n293 ? n441 : !n441)));
assign n820  = /* LUT    8 12  1 */ (n371 ? (n433 ? (n188 ? 1'b1 : n455) : 1'b1) : (n433 ? 1'b1 : (n188 ? n455 : 1'b1)));
assign n821  = /* LUT    2 12  7 */ n55;
assign n822  = /* LUT    9  5  5 */ n471;
assign n823  = /* LUT    6  4  4 */ n218;
assign n824  = /* LUT    6  7  6 */ n237;
assign n825  = /* LUT    9  6  6 */ (n107 ? (n7 ? n485 : n477) : n485);
assign n826  = /* LUT    7  9  0 */ (n10 ? (n337 ? n168 : !n168) : (n337 ? !n168 : n168));
assign n827  = /* LUT   11 11  5 */ n529;
assign n828  = /* LUT   11  3  1 */ (n313 ? (n209 ? !n444 : n444) : (n209 ? n444 : !n444));
assign n829  = /* LUT    6 11  3 */ (n270 ? (n38 ? 1'b1 : (n58 ? 1'b1 : n52)) : 1'b0);
assign n830  = /* LUT    8 11  5 */ (n416 ? !n348 : n348);
assign n831  = /* LUT    7 12  1 */ (n351 ? (n367 ? !n441 : n441) : (n367 ? n441 : !n441));
assign n832  = /* LUT    2  8  5 */ (n32 ? (n42 ? n20 : n22) : (n42 ? !n20 : !n22));
assign n833  = /* LUT    5  4  4 */ (n146 ? (n8 ? n83 : !n83) : (n8 ? !n83 : n83));
assign n834  = /* LUT    6  8  6 */ (n42 ? n247 : n256);
assign n835  = /* LUT    4  8  7 */ n32;
assign n836  = /* LUT    7  4  6 */ (n101 ? n297 : !n112);
assign n837  = /* LUT    7 13  2 */ (n133 ? !n280 : n280);
assign n838  = /* LUT    5  5  5 */ n148;
assign n839  = /* LUT    9  5  0 */ n468;
assign n840  = /* LUT    2 12  2 */ n57;
assign n841  = /* LUT    7  5  7 */ n311;
assign n842  = /* LUT    4 12  4 */ (n117 ? 1'b0 : !n116);
assign n843  = /* LUT    6  7  1 */ (n107 ? (n7 ? n102 : 1'b1) : (n7 ? n240 : 1'b0));
assign n844  = /* LUT    8  7  3 */ (n407 ? (n167 ? (n403 ? !n15 : 1'b1) : (n403 ? n15 : 1'b0)) : (n167 ? (n403 ? n15 : 1'b0) : (n403 ? !n15 : 1'b1)));
assign n845  = /* LUT    5  8  6 */ n171;
assign n846  = /* LUT    9  8  1 */ n487;
assign n847  = /* LUT    4 15  5 */ (n52 ? !n131 : 1'b0);
assign n848  = /* LUT    7 11  4 */ (n336 ? (n353 ? !n201 : 1'b0) : (n353 ? n352 : 1'b1));
assign n849  = /* LUT    4  7  1 */ n44;
assign n850  = /* LUT    8 11  0 */ (n421 ? (n506 ? (n347 ? n344 : !n344) : n347) : (n506 ? 1'b1 : n344));
assign n851  = /* LUT    6 11  7 */ n257;
assign n852  = /* LUT   11  6  7 */ n518;
assign n853  = /* LUT   11  9  3 */ n257;
assign n854  = /* LUT    5 12  3 */ (n192 ? (n196 ? 1'b0 : !n193) : (n196 ? !n191 : (n193 ? !n191 : n191)));
assign n855  = /* LUT    7 12  5 */ (n2 ? (n433 ? (n188 ? n437 : 1'b0) : 1'b0) : 1'b0);
assign n856  = /* LUT    6  8  1 */ (n106 ? (n15 ? n247 : 1'b0) : (n15 ? !n247 : 1'b1));
assign n857  = /* LUT    4  8  2 */ n100;
assign n858  = /* LUT    7  4  1 */ (n107 ? (n7 ? !n297 : 1'b1) : (n7 ? !n302 : 1'b0));
assign n859  = /* LUT    8  8  3 */ n404;
assign n860  = /* LUT   11 10  4 */ !n529;
assign n861  = /* LUT    5  5  0 */ n151;
assign n862  = /* LUT    7  5  2 */ (n7 ? (n107 ? n309 : n226) : n309);
assign n863  = /* LUT    9  5  4 */ n466;
assign n864  = /* LUT    2  4  2 */ n12;
assign n865  = /* LUT    4 11  3 */ n28;
assign n866  = /* LUT    6 15  0 */ (n286 ? (n274 ? !n285 : n285) : 1'b0);
assign n867  = /* LUT    6  7  5 */ n239;
assign n868  = /* LUT    8  7  7 */ (n167 ? (n15 ? !n72 : 1'b1) : (n15 ? n72 : 1'b0));
assign n869  = /* LUT   11 13  5 */ (n542 ? !n188 : n188);
assign n870  = /* LUT    5  8  1 */ n174;
assign n871  = /* LUT    4 15  0 */ (n38 ? (n63 ? (n205 ? n129 : 1'b1) : 1'b0) : (n205 ? n129 : 1'b1));
assign n872  = /* LUT    9  8  5 */ n489;
assign n873  = /* LUT    5 11  6 */ (n263 ? !n202 : n202);
assign n874  = /* LUT    2  7  3 */ n16;
assign n875  = /* LUT    4  7  5 */ n85;
assign n876  = /* LUT    6 11  2 */ (n192 ? (n30 ? 1'b1 : n266) : (n30 ? n191 : (n266 ? n191 : !n191)));
assign n877  = /* LUT    8 11  4 */ (n421 ? (n506 ? !n344 : (n347 ? !n344 : n344)) : (n506 ? 1'b0 : !n347));
assign n878  = /* LUT   11  9  7 */ (n209 ? (n15 ? n525 : 1'b0) : (n15 ? !n525 : 1'b1));
assign n879  = /* LUT    7 12  0 */ (n2 ? !n439 : 1'b0);
assign n880  = /* LUT    5  4  3 */ (n11 ? (n6 ? n189 : 1'b1) : (n6 ? !n189 : 1'b0));
assign n881  = /* LUT    4  8  6 */ n95;
assign n882  = /* LUT    7  4  5 */ (n7 ? (n107 ? n302 : n297) : n302);
assign n883  = /* LUT    6  3  3 */ (n10 ? (n15 ? !n215 : 1'b1) : (n15 ? n215 : 1'b0));
assign n884  = /* LUT    8 14  5 */ (n357 ? (n278 ? n451 : 1'b1) : (n452 ? (n278 ? 1'b1 : n451) : (n278 ? 1'b0 : !n451)));
assign n885  = /* LUT    7 15  1 */ (n286 ? (n374 ? 1'b0 : (n363 ? n290 : 1'b1)) : 1'b0);
assign n886  = /* LUT    5  7  4 */ (n242 ? (n15 ? n71 : 1'b0) : (n15 ? !n71 : 1'b1));
assign n887  = /* LUT    6 15  4 */ (n189 ? !n52 : 1'b0);
assign n888  = /* LUT    7  7  6 */ n325;
assign n889  = /* LUT    4  3  3 */ n82;
assign n890  = /* LUT    6  7  0 */ (n235 ? (n7 ? 1'b1 : n161) : (n7 ? 1'b0 : !n48));
assign n891  = /* LUT    4 14  3 */ (n207 ? (n125 ? 1'b0 : !n130) : (n125 ? !n130 : 1'b0));
assign n892  = /* LUT    8  7  2 */ (n167 ? (n15 ? !n50 : 1'b1) : (n15 ? n50 : 1'b0));
assign n896  = /* LUT   11  5  5 */ n514;
assign n897  = /* LUT    5  8  5 */ (n106 ? (n168 ? (n21 ? n15 : 1'b0) : (n21 ? !n15 : 1'b1)) : (n168 ? (n21 ? !n15 : 1'b1) : (n21 ? n15 : 1'b0)));
assign n898  = /* LUT    9  8  0 */ n500;
assign n899  = /* LUT    2 15  2 */ (rst ? 1'b0 : (n64 ? 1'b1 : (n38 ? n63 : 1'b0)));
assign n900  = /* LUT    5 11  1 */ (n163 ? (n38 ? 1'b0 : (n58 ? 1'b0 : !n52)) : 1'b0);
assign n901  = /* LUT    4 15  4 */ (n127 ? (n126 ? (n124 ? !n125 : 1'b0) : 1'b0) : 1'b0);
assign n902  = /* LUT    7 11  3 */ (n336 ? (n201 ? (n352 ? 1'b0 : !n353) : n352) : (n201 ? (n352 ? 1'b0 : n353) : 1'b1));
assign n903  = /* LUT    4  7  0 */ n87;
assign n904  = /* LUT    2  7  7 */ (n42 ? n71 : n45);
assign n905  = /* LUT   11  6  6 */ n165;
assign n906  = /* LUT   11  9  2 */ (n42 ? n526 : n523);
assign n907  = /* LUT    7 12  4 */ (n2 ? !n434 : 1'b0);
assign n908  = /* LUT    4  8  1 */ n94;
assign n909  = /* LUT    7  4  0 */ (n300 ? (n7 ? 1'b1 : !n306) : (n7 ? 1'b0 : n112));
assign n910  = /* LUT    8 14  0 */ (n363 ? (n208 ? (n362 ? 1'b0 : n132) : n362) : (n208 ? (n362 ? 1'b0 : !n132) : 1'b1));
assign n911  = /* LUT    8  3  0 */ (n378 ? (n7 ? 1'b1 : !n379) : (n7 ? 1'b0 : n65));
assign n912  = /* LUT    6  3  7 */ (n10 ? (n15 ? !n213 : 1'b1) : (n15 ? n213 : 1'b0));
assign n913  = /* LUT    6 14  7 */ (n279 ? (n288 ? (n36 ? 1'b1 : n357) : (n36 ? 1'b0 : !n357)) : (n288 ? (n36 ? 1'b0 : !n357) : (n36 ? 1'b1 : n357)));
assign n914  = /* LUT    4 11  2 */ (n38 ? 1'b0 : (n58 ? 1'b0 : !n52));
assign n915  = /* LUT    7  7  1 */ (n107 ? (n7 ? n314 : 1'b1) : (n7 ? n328 : 1'b0));
assign n916  = /* LUT    9  4  7 */ n464;
assign n917  = /* LUT    9  7  3 */ (n107 ? (n7 ? n332 : n248) : n332);
assign n918  = /* LUT    4  3  7 */ n79;
assign n919  = /* LUT    6  7  4 */ (n101 ? n102 : !n48);
assign n920  = /* LUT    8  7  6 */ n400;
assign n921  = /* LUT   11 13  4 */ (n541 ? !n433 : n433);
assign n922  = /* LUT   11  5  0 */ (n107 ? 1'b0 : !n7);
assign n923  = /* LUT    5  8  0 */ n96;
assign n924  = /* LUT    9  8  4 */ n488;
assign n925  = /* LUT    2 15  6 */ (rst ? 1'b0 : (n58 ? 1'b1 : (n38 ? !n63 : 1'b0)));
assign n926  = /* LUT    2  7  2 */ n17;
assign n927  = /* LUT   11  6  1 */ n29;
assign n928  = /* LUT    5 14  7 */ (n205 ? 1'b0 : (n38 ? 1'b0 : (n58 ? 1'b0 : !n2)));
assign n929  = /* LUT    6 10  5 */ (n259 ? (n263 ? (n202 ? 1'b1 : n189) : (n202 ? n189 : 1'b1)) : (n263 ? (n202 ? 1'b0 : !n189) : (n202 ? !n189 : 1'b0)));
assign n930  = /* LUT   11  9  6 */ (n406 ? (n209 ? (n528 ? !n15 : 1'b1) : (n528 ? n15 : 1'b0)) : (n209 ? (n528 ? n15 : 1'b0) : (n528 ? !n15 : 1'b1)));
assign n931  = /* LUT    8 10  7 */ (n397 ? (n416 ? (n498 ? n422 : 1'b1) : (n498 ? !n422 : 1'b0)) : (n498 ? !n422 : 1'b0));
assign n932  = /* LUT    9 11  5 */ (n502 ? (n510 ? !n509 : n509) : (n510 ? n509 : !n509));
assign n933  = /* LUT    5  3  6 */ n140;
assign n934  = /* LUT    4 10  5 */ n104;
assign n935  = /* LUT    6 14  2 */ (n273 ? (n278 ? n277 : !n277) : (n278 ? !n277 : n277));
assign n936  = /* LUT    6  3  2 */ (n42 ? n215 : n210);
assign n937  = /* LUT    8 14  4 */ (n36 ? (n77 ? 1'b1 : n452) : (n77 ? n451 : (n452 ? n451 : !n451)));
assign n938  = /* LUT    8  3  4 */ n382;
assign n939  = /* LUT    7 15  0 */ (n292 ? n453 : !n453);
assign n940  = /* LUT   11  4  3 */ (n313 ? !n444 : n444);
assign n941  = /* LUT    5 15  7 */ (rst ? 1'b0 : (n2 ? 1'b1 : (n205 ? !n129 : 1'b0)));
assign n942  = /* LUT    5  7  3 */ n19;
assign n943  = /* LUT    4 11  6 */ n183;
assign n944  = /* LUT    7  7  5 */ n329;
assign n945  = /* LUT    4  3  2 */ n80;
assign n946  = /* LUT    4 14  2 */ (n206 ? (n124 ? 1'b0 : !n130) : (n124 ? !n130 : 1'b0));
assign n947  = /* LUT    9  7  7 */ n495;
assign n948  = /* LUT    8  7  1 */ (n407 ? (n15 ? n405 : 1'b0) : (n15 ? !n405 : 1'b1));
assign n949  = /* LUT    8  6  5 */ (n53 ? !n88 : n88);
assign n950  = /* LUT    5 11  0 */ (n110 ? (n38 ? 1'b1 : (n58 ? 1'b1 : n52)) : 1'b0);
assign n951  = /* LUT    7 11  2 */ (n352 ? (n336 ? (n353 ? !n201 : n201) : (n353 ? n201 : 1'b0)) : (n336 ? (n353 ? 1'b0 : !n201) : 1'b1));
assign n952  = /* LUT    7 14  4 */ (n372 ? (n133 ? !n369 : 1'b1) : (n133 ? n369 : 1'b0));
assign n953  = /* LUT    6 10  0 */ n254;
assign n954  = /* LUT   11  9  1 */ (n42 ? n527 : n537);
assign n955  = /* LUT    8 10  2 */ (n415 ? !n334 : n334);
assign n956  = /* LUT    6 13  5 */ (n269 ? (n74 ? !n198 : n198) : (n74 ? n198 : !n198));
assign n957  = /* LUT    9 11  0 */ (n507 ? (n416 ? (n348 ? 1'b0 : !n421) : (n348 ? !n421 : 1'b0)) : (n416 ? (n348 ? 1'b1 : n421) : (n348 ? n421 : 1'b1)));
assign n958  = /* LUT    5  3  1 */ n40;
assign n959  = /* LUT    7  3  3 */ n299;
assign n960  = /* LUT    9  3  5 */ n458;
assign n961  = /* LUT    5  6  6 */ (n209 ? (n15 ? n156 : 1'b0) : (n15 ? !n156 : 1'b1));
assign n962  = /* LUT    6 14  6 */ (n278 ? !n77 : 1'b0);
assign n963  = /* LUT    6  6  2 */ n233;
assign n964  = /* LUT    5 15  2 */ (rst ? 1'b0 : !n62);
assign n965  = /* LUT    7 15  4 */ (n291 ? n453 : !n453);
assign n966  = /* LUT    7  7  0 */ (n323 ? (n7 ? 1'b0 : !n331) : (n7 ? 1'b1 : n103));
assign n967  = /* LUT    9  4  6 */ n462;
assign n968  = /* LUT    5  7  7 */ n164;
assign n969  = /* LUT    9  7  2 */ (n479 ? (n7 ? 1'b1 : !n332) : (n7 ? 1'b0 : n492));
assign n970  = /* LUT   11 13  3 */ (n540 ? !n534 : n534);
assign n971  = /* LUT    6  9  3 */ (n8 ? (n15 ? !n251 : 1'b1) : (n15 ? n251 : 1'b0));
assign n972  = /* LUT    8  9  5 */ (n341 ? (n420 ? (n428 ? n338 : !n338) : (n428 ? !n338 : n338)) : (n420 ? (n428 ? !n338 : n338) : (n428 ? n338 : !n338)));
assign n973  = /* LUT    9 14  1 */ (rst ? 1'b1 : (n123 ? !n39 : 1'b0));
assign n974  = /* LUT    4  6  7 */ n6;
assign n975  = /* LUT    6 10  4 */ n26;
assign n976  = /* LUT    6 13  0 */ (n75 ? !n198 : n198);
assign n977  = /* LUT    8 10  6 */ (n432 ? (n497 ? (n498 ? !n431 : n431) : !n498) : (n497 ? !n431 : 1'b0));
assign n978  = /* LUT    9 11  4 */ (n511 ? (n504 ? !n501 : n501) : (n504 ? n501 : !n501));
assign n979  = /* LUT    5  3  5 */ n184;
assign n980  = /* LUT    5  6  1 */ (n209 ? (n15 ? n157 : 1'b0) : (n15 ? !n157 : 1'b1));
assign n981  = /* LUT    8 14  3 */ (n77 ? (n36 ? 1'b0 : (n278 ? n357 : !n357)) : (n36 ? (n278 ? n357 : !n357) : 1'b0));
assign n982  = /* LUT    8 13  7 */ (n356 ? (n445 ? (n433 ? 1'b0 : !n371) : 1'b1) : (n445 ? (n433 ? 1'b1 : n371) : 1'b0));
assign n983  = /* LUT    9  4  1 */ n461;
assign n984  = /* LUT    5  7  2 */ (n242 ? (n15 ? n70 : 1'b0) : (n15 ? !n70 : 1'b1));
assign n985  = /* LUT    7  7  4 */ (n101 ? n314 : !n103);
assign n986  = /* LUT    4  3  1 */ (n10 ? !n6 : n6);
assign n989  = /* LUT    9  7  6 */ n483;
assign n990  = /* LUT    5 10  4 */ n163;
assign n991  = /* LUT    7 10  6 */ (n339 ? (n340 ? (n427 ? !n418 : n418) : (n427 ? n418 : !n418)) : (n340 ? (n427 ? n418 : !n418) : (n427 ? !n418 : n418)));
assign n992  = /* LUT    8  6  4 */ (n101 ? n392 : !n47);
assign n993  = /* LUT    8  9  0 */ (n397 ? (n307 ? (n377 ? n159 : !n159) : (n377 ? !n159 : n159)) : (n307 ? (n377 ? !n159 : n159) : (n377 ? n159 : !n159)));
assign n994  = /* LUT    6  9  7 */ n253;
assign n995  = /* LUT    7 14  3 */ (n375 ? (n293 ? (n369 ? n285 : 1'b1) : (n369 ? !n285 : 1'b0)) : (n293 ? (n369 ? !n285 : 1'b0) : (n369 ? n285 : 1'b1)));
assign n996  = /* LUT    8 10  1 */ (n415 ? (n496 ? !n334 : n334) : (n496 ? n334 : !n334));
assign n997  = /* LUT    6 13  4 */ (n277 ? (n269 ? (n122 ? !n276 : n276) : !n276) : (n269 ? 1'b1 : !n122));
assign n998  = /* LUT    7  3  2 */ (n107 ? (n7 ? n306 : n297) : n306);
assign n999  = /* LUT    9  3  4 */ (n107 ? (n7 ? n379 : n460) : n379);
assign n1000 = /* LUT    2 10  6 */ n54;
assign n1001 = /* LUT    5  6  5 */ (n166 ? (n209 ? (n14 ? !n15 : 1'b1) : (n14 ? n15 : 1'b0)) : (n209 ? (n14 ? n15 : 1'b0) : (n14 ? !n15 : 1'b1)));
assign n1002 = /* LUT    7  6  4 */ (n107 ? (n7 ? n331 : n314) : n331);
assign n1003 = /* LUT   11 12  1 */ (n371 ? (n433 ? (n455 ? 1'b0 : !n188) : 1'b0) : 1'b0);
assign n1004 = /* LUT    8 13  2 */ (n35 ? (n442 ? (n448 ? !n360 : n360) : (n448 ? n360 : !n360)) : 1'b0);
assign n1005 = /* LUT    5  9  7 */ (n166 ? (n178 ? !n15 : 1'b1) : (n178 ? n15 : 1'b0));
assign n1006 = /* LUT    1 12  0 */ n33;
assign n1007 = /* LUT    6  5  5 */ n223;
assign n1008 = /* LUT    8  5  7 */ n393;
assign n1009 = /* LUT    7 10  1 */ (n424 ? !n427 : n427);
assign n1010 = /* LUT    9 10  3 */ (n478 ? (n264 ? n334 : !n334) : (n264 ? !n334 : n334));
assign n1011 = /* LUT    6  9  2 */ (n242 ? (n15 ? n243 : 1'b0) : (n15 ? !n243 : 1'b1));
assign n1012 = /* LUT    8  9  4 */ (n425 ? n418 : !n418);
assign n1013 = /* LUT   11  7  7 */ (n42 ? n50 : n522);
assign n1014 = /* LUT    2  6  4 */ n14;
assign n1015 = /* LUT   12  7  3 */ n536;
assign n1016 = /* LUT    7 14  7 */ (n208 ? (n132 ? (n363 ? 1'b1 : n362) : (n363 ? n362 : 1'b1)) : (n132 ? 1'b0 : n362));
assign n1017 = /* LUT    6 12  3 */ (n232 ? (n283 ? (n354 ? 1'b1 : !n35) : (n354 ? !n35 : 1'b1)) : (n283 ? (n354 ? 1'b0 : n35) : (n354 ? n35 : 1'b0)));
assign n1018 = /* LUT    8 12  5 */ (n455 ? !n371 : (n188 ? !n371 : n433));
assign n1019 = /* LUT    5  6  0 */ (n104 ? (n42 ? n154 : n158) : (n42 ? !n154 : !n158));
assign n1020 = /* LUT    9  6  1 */ n474;
assign n1021 = /* LUT    5  9  2 */ (n53 ? (n15 ? !n179 : 1'b1) : (n15 ? n179 : 1'b0));
assign n1022 = /* LUT    7  9  4 */ (n340 ? (n418 ? (n255 ? !n15 : 1'b1) : (n255 ? n15 : 1'b0)) : (n418 ? (n255 ? n15 : 1'b0) : (n255 ? !n15 : 1'b1)));
assign n1023 = /* LUT    6  5  0 */ n217;
assign n1024 = /* LUT    8 13  6 */ (n454 ? (n358 ? (n450 ? n364 : !n364) : (n450 ? !n364 : n364)) : (n358 ? (n450 ? !n364 : n364) : (n450 ? n364 : !n364)));
assign n1025 = /* LUT   11 11  0 */ (n76 ? n34 : 1'b0);
assign n1026 = /* LUT    9  9  6 */ n187;
assign n1027 = /* LUT    8  5  2 */ n395;
assign n1028 = /* LUT    7 10  5 */ (n264 ? (n346 ? (n343 ? !n423 : n423) : !n343) : (n346 ? n423 : 1'b0));
assign n1029 = /* LUT    9 10  7 */ (n264 ? !n159 : 1'b0);
assign n1030 = /* LUT    6  9  6 */ n335;
assign n1031 = /* LUT    4  9  7 */ n178;
assign n1032 = /* LUT   11  7  2 */ n481;
assign n1033 = /* LUT    4  6  1 */ (n160 ? !n84 : n84);
assign n1034 = /* LUT    7 14  2 */ (n132 ? (n208 ? (n362 ? 1'b1 : n363) : (n362 ? n363 : 1'b1)) : (n208 ? 1'b0 : n363));
assign n1035 = /* LUT    7 13  6 */ (n358 ? (n368 ? (n450 ? !n364 : n364) : (n450 ? n364 : !n364)) : (n368 ? (n450 ? n364 : !n364) : (n450 ? !n364 : n364)));
assign n1036 = /* LUT   11  8  3 */ n403;
assign n1037 = /* LUT    8 12  0 */ (n412 ? (n440 ? (n443 ? 1'b1 : !n35) : (n443 ? !n35 : 1'b1)) : (n440 ? (n443 ? 1'b0 : n35) : (n443 ? n35 : 1'b0)));
assign n1038 = /* LUT    2 12  6 */ n61;
assign n1039 = /* LUT    6 12  7 */ (n192 ? 1'b0 : !n191);
assign n1040 = /* LUT    6  4  3 */ n219;
assign n1041 = /* LUT    8  4  5 */ n386;
assign n1042 = /* LUT    7  6  3 */ n319;
assign n1043 = /* LUT    9  6  5 */ n104;
assign n1044 = /* LUT    2 13  7 */ (n38 ? 1'b0 : !n52);
assign n1045 = /* LUT    5  9  6 */ (n42 ? n179 : n180);
assign n1046 = /* LUT    8 13  1 */ (n355 ? (n446 ? !n441 : n441) : (n446 ? n441 : !n441));
assign n1047 = /* LUT    9  9  1 */ (n499 ? !n478 : n478);
assign n1048 = /* LUT    6  5  4 */ n228;
assign n1049 = /* LUT    8  5  6 */ (n7 ? (n107 ? n391 : n392) : n391);
assign n1050 = /* LUT   11 11  4 */ (n76 ? 1'b1 : (n530 ? (n534 ? 1'b1 : n34) : 1'b0));
assign n1051 = /* LUT    9 10  2 */ (n498 ? (n503 ? 1'b0 : (n506 ? n421 : !n421)) : (n503 ? (n506 ? n421 : !n421) : 1'b0));
assign n1052 = /* LUT    8  9  3 */ (n419 ? (n338 ? (n425 ? !n418 : n418) : (n425 ? n418 : !n418)) : (n338 ? (n425 ? n418 : !n418) : (n425 ? !n418 : n418)));
assign n1053 = /* LUT   11  7  6 */ n520;
assign n1054 = /* LUT    8  8  7 */ n408;
assign n1055 = /* LUT    7 13  1 */ (n122 ? (n365 ? !n277 : 1'b0) : (n365 ? (n277 ? n370 : !n370) : !n370));
assign n1056 = /* LUT    9 13  3 */ !n76;
assign n1057 = /* LUT    2 12  1 */ (n57 ? (n38 ? 1'b0 : (n58 ? 1'b0 : !n52)) : 1'b0);
assign n1058 = /* LUT    7  5  6 */ (n101 ? n226 : !n229);
assign n1059 = /* LUT    6 12  2 */ (n267 ? (n190 ? 1'b1 : n197) : (n190 ? 1'b0 : !n197));
assign n1060 = /* LUT    4 12  3 */ (n120 ? (n38 ? 1'b1 : (n58 ? 1'b1 : n52)) : 1'b0);
assign n1061 = /* LUT    8 12  4 */ (n455 ? !n371 : 1'b0);
assign n1062 = /* LUT    8  4  0 */ n388;
assign n1063 = /* LUT    6  4  7 */ (n160 ? (n167 ? n84 : !n84) : (n167 ? !n84 : n84));
assign n1064 = /* LUT    9  6  0 */ (n107 ? (n7 ? !n477 : 1'b1) : (n7 ? 1'b1 : n402));
assign n1065 = /* LUT    5  9  1 */ (n176 ? (n42 ? n177 : n181) : (n42 ? !n177 : !n181));
assign n1066 = /* LUT    7  6  7 */ n316;
assign n1067 = /* LUT    7  9  3 */ (n10 ? !n337 : n337);
assign n1068 = /* LUT    8 13  5 */ (n449 ? !n280 : 1'b0);
assign n1069 = /* LUT    9  9  5 */ (n480 ? !n377 : n377);
assign n1070 = /* LUT    8  5  1 */ n401;
assign n1071 = /* LUT    6 11  6 */ (n254 ? (n38 ? 1'b0 : (n58 ? 1'b0 : !n52)) : 1'b0);
assign n1072 = /* LUT    6  8  0 */ n176;
assign n1073 = /* LUT    8  8  2 */ n414;
assign n1074 = /* LUT    5  4  7 */ n144;
assign n1075 = /* LUT    7 13  5 */ (n359 ? !n293 : n293);
assign n1076 = /* LUT    7  5  1 */ (n107 ? (n7 ? !n226 : 1'b1) : (n7 ? !n309 : 1'b0));
assign n1077 = /* LUT   12  9  6 */ n528;
assign n1078 = /* LUT    9  5  3 */ n470;
assign n1079 = /* LUT    6 12  6 */ (n272 ? (n75 ? (n267 ? !n199 : n199) : (n267 ? n199 : !n199)) : (n75 ? (n267 ? n199 : !n199) : (n267 ? !n199 : n199)));
assign n1080 = /* LUT    4 12  7 */ n32;
assign n1081 = /* LUT    6  4  2 */ n142;
assign n1082 = /* LUT    8  4  4 */ n380;
assign n1083 = /* LUT    7  6  2 */ n320;
assign n1084 = /* LUT    9  6  4 */ (n101 ? n477 : !n402);
assign n1085 = /* LUT    5  9  5 */ (n42 ? n182 : n105);
assign n1086 = /* LUT    9  9  0 */ (n480 ? n397 : !n397);
assign n1087 = /* LUT    2  5  2 */ n41;
assign n1088 = /* LUT    7  9  7 */ (n409 ? !n321 : n321);
assign n1089 = /* LUT    6 11  1 */ (n29 ? (n38 ? 1'b0 : (n58 ? 1'b0 : !n52)) : 1'b0);
assign n1090 = /* LUT    8 11  3 */ (n159 ? !n497 : n497);
assign n540  = /* CARRY 11 13  2 */ (1'b0 & n530) | ((1'b0 | n530) & n539);
assign n545  = /* CARRY  4 14  0 */ (n127 & 1'b0) | ((n127 | 1'b0) & n664);
assign n544  = /* CARRY 11 13  6 */ (1'b0 & n455) | ((1'b0 | n455) & n543);
assign n539  = /* CARRY 11 13  1 */ (1'b0 & n34) | ((1'b0 | n34) & n546);
assign n543  = /* CARRY 11 13  5 */ (1'b0 & n188) | ((1'b0 | n188) & n542);
assign n546  = /* CARRY 11 13  0 */ (n76 & 1'b0) | ((n76 | 1'b0) & n895);
assign n542  = /* CARRY 11 13  4 */ (1'b0 & n433) | ((1'b0 | n433) & n541);
assign n207  = /* CARRY  4 14  2 */ (1'b0 & n124) | ((1'b0 | n124) & n206);
assign n541  = /* CARRY 11 13  3 */ (1'b0 & n534) | ((1'b0 | n534) & n540);
assign n206  = /* CARRY  4 14  1 */ (1'b0 & n126) | ((1'b0 | n126) & n545);
/* FF  5 12  6 */ always @(posedge clk) if (n2) n200 <= 1'b0 ? 1'b0 : n547;
/* FF  9 12  1 */ assign n203 = n548;
/* FF  5  4  2 */ always @(posedge clk) if (1'b1) n142 <= 1'b0 ? 1'b0 : n549;
/* FF  4  8  5 */ always @(posedge clk) if (1'b1) n99 <= 1'b0 ? 1'b0 : n550;
/* FF  8  8  6 */ always @(posedge clk) if (1'b1) n413 <= 1'b0 ? 1'b0 : n551;
/* FF  7  4  4 */ always @(posedge clk) if (1'b1) n303 <= 1'b0 ? 1'b0 : n552;
/* FF  7 13  0 */ assign n355 = n553;
/* FF  9 13  2 */ assign n513 = n554;
/* FF  5  5  3 */ always @(posedge clk) if (1'b1) n150 <= 1'b0 ? 1'b0 : n555;
/* FF  6 12  1 */ assign n272 = n556;
/* FF  7  5  5 */ always @(posedge clk) if (1'b1) n310 <= 1'b0 ? 1'b0 : n557;
/* FF  4 12  2 */ assign n117 = n558;
/* FF  8 12  3 */ assign n436 = n559;
/* FF  6 15  3 */ assign n291 = n560;
/* FF  5  9  0 */ assign n166 = n561;
/* FF  9  9  4 */ assign n498 = n562;
/* FF  5  8  4 */ always @(posedge clk) if (1'b1) n174 <= 1'b0 ? 1'b0 : n563;
/* FF  7  8  6 */ always @(posedge clk) if (1'b1) n255 <= 1'b0 ? 1'b0 : n564;
/* FF  4 15  3 */ assign n130 = n565;
/* FF 11  6  5 */ always @(posedge clk) if (1'b1) n517 <= 1'b0 ? 1'b0 : n566;
/* FF  8 11  7 */ assign n432 = n567;
/* FF  5 12  1 */ assign n197 = n568;
/* FF  7 12  3 */ assign n84 = n569;
/* FF  4  8  0 */ always @(posedge clk) if (1'b1) n94 <= 1'b0 ? 1'b0 : n570;
/* FF  8  8  1 */ always @(posedge clk) if (1'b1) n408 <= 1'b0 ? 1'b0 : n571;
/* FF  5  4  6 */ always @(posedge clk) if (1'b1) n145 <= 1'b0 ? 1'b0 : n572;
/* FF  7 13  4 */ assign n359 = n573;
/* FF  7  5  0 */ assign n307 = n574;
/* FF  5  5  7 */ always @(posedge clk) if (1'b1) n153 <= 1'b0 ? 1'b0 : n575;
/* FF  9  5  2 */ always @(posedge clk) if (1'b1) n467 <= 1'b0 ? 1'b0 : n576;
/* FF  2 12  4 */ always @(posedge clk) if (1'b1) n55 <= 1'b0 ? 1'b0 : n577;
/* FF  2  4  0 */ always @(posedge clk) if (1'b1) n41 <= 1'b0 ? 1'b0 : n578;
/* FF  4 12  6 */ always @(posedge clk) if (n2) n119 <= 1'b0 ? 1'b0 : n579;
/* FF  6 15  7 */ assign n292 = n580;
/* FF  6  7  3 */ always @(posedge clk) if (1'b1) n236 <= 1'b0 ? 1'b0 : n581;
/* FF  7  8  1 */ always @(posedge clk) if (1'b1) n330 <= 1'b0 ? 1'b0 : n582;
/* FF  5 11  4 */ assign n193 = n583;
/* FF  4 15  7 */ assign n62 = n584;
/* FF  7 11  6 */ assign n347 = n585;
/* FF  4  7  3 */ always @(posedge clk) if (1'b1) n91 <= 1'b0 ? 1'b0 : n586;
/* FF 11  6  0 */ assign n493 = n587;
/* FF  8 11  2 */ assign n427 = n588;
/* FF 11  9  5 */ always @(posedge clk) if (1'b1) n526 <= 1'b0 ? 1'b0 : n589;
/* FF  5 12  5 */ assign n33 = n590;
/* FF  7 12  7 */ assign n351 = n591;
/* FF  5  4  1 */ always @(posedge clk) if (1'b1) n9 <= 1'b0 ? 1'b0 : n592;
/* FF  6  8  3 */ always @(posedge clk) if (1'b1) n22 <= 1'b0 ? 1'b0 : n593;
/* FF  4  8  4 */ always @(posedge clk) if (1'b1) \d_out[7]  <= 1'b0 ? 1'b0 : n594;
/* FF  7  4  3 */ always @(posedge clk) if (1'b1) n302 <= 1'b0 ? 1'b0 : n595;
/* FF  8  8  5 */ always @(posedge clk) if (1'b1) n412 <= 1'b0 ? 1'b0 : n596;
/* FF  6  3  1 */ always @(posedge clk) if (1'b1) n211 <= 1'b0 ? 1'b0 : n597;
/* FF  6 14  1 */ assign n285 = n598;
/* FF  8  3  3 */ always @(posedge clk) if (1'b1) n380 <= 1'b0 ? 1'b0 : n599;
/* FF  6  6  6 */ always @(posedge clk) if (1'b1) n233 <= 1'b0 ? 1'b0 : n600;
/* FF  4 11  5 */ always @(posedge clk) if (1'b1) n59 <= 1'b0 ? 1'b0 : n601;
/* FF  6 15  2 */ assign n290 = n602;
/* FF  8  7  0 */ assign n402 = n603;
/* FF  6  7  7 */ always @(posedge clk) if (1'b1) n240 <= 1'b0 ? 1'b0 : n604;
/* FF 11 13  7 */ always @(posedge clk) if (1'b1) n371 <= n3 ? 1'b0 : n605;
/* FF  5  8  3 */ always @(posedge clk) if (1'b1) n173 <= 1'b0 ? 1'b0 : n606;
/* FF  7  8  5 */ always @(posedge clk) if (1'b1) n331 <= 1'b0 ? 1'b0 : n607;
/* FF  4 15  2 */ assign n129 = n608;
/* FF  9  8  7 */ always @(posedge clk) if (1'b1) n23 <= 1'b0 ? 1'b0 : n609;
/* FF  7 11  1 */ assign n343 = n610;
/* FF  4  7  7 */ always @(posedge clk) if (1'b1) n93 <= 1'b0 ? 1'b0 : n611;
/* FF  6 11  4 */ assign n269 = n612;
/* FF  8 11  6 */ assign n431 = n613;
/* FF 11  6  4 */ always @(posedge clk) if (1'b1) n485 <= 1'b0 ? 1'b0 : n614;
/* FF 11  9  0 */ assign n492 = n615;
/* FF  5 12  0 */ assign n196 = n616;
/* FF  7 12  2 */ assign n202 = n617;
/* FF  5  4  5 */ always @(posedge clk) if (1'b1) n144 <= 1'b0 ? 1'b0 : n618;
/* FF  2 11  2 */ assign n30 = n619;
/* FF  7  4  7 */ always @(posedge clk) if (1'b1) n306 <= 1'b0 ? 1'b0 : n620;
/* FF  6  3  5 */ always @(posedge clk) if (1'b1) n215 <= 1'b0 ? 1'b0 : n621;
/* FF  6 14  5 */ assign n287 = n622;
/* FF  8 14  7 */ assign n293 = n623;
/* FF  6  6  1 */ assign n229 = n624;
/* FF  8  3  7 */ always @(posedge clk) if (1'b1) n383 <= 1'b0 ? 1'b0 : n625;
/* FF  4 11  0 */ assign n113 = n626;
/* FF  5  7  6 */ always @(posedge clk) if (1'b1) n164 <= 1'b0 ? 1'b0 : n627;
/* FF  9  7  1 */ assign n479 = n628;
/* FF  2  3  3 */ always @(posedge clk) if (1'b1) n40 <= 1'b0 ? 1'b0 : n629;
/* FF  4 14  5 */ always @(posedge clk) if (n121) n127 <= rst ? 1'b0 : n630;
/* FF  6  7  2 */ always @(posedge clk) if (1'b1) n16 <= 1'b0 ? 1'b0 : n631;
/* FF 11 13  2 */ always @(posedge clk) if (1'b1) n530 <= n3 ? 1'b0 : n632;
/* FF  5  8  7 */ always @(posedge clk) if (1'b1) n21 <= 1'b0 ? 1'b0 : n633;
/* FF  9  8  2 */ always @(posedge clk) if (1'b1) n489 <= 1'b0 ? 1'b0 : n634;
/* FF  5 11  3 */ assign n192 = n635;
/* FF  2  7  0 */ always @(posedge clk) if (1'b1) n45 <= 1'b0 ? 1'b0 : n636;
/* FF  4 15  6 */ assign n131 = n637;
/* FF  4  7  2 */ always @(posedge clk) if (1'b1) n67 <= 1'b0 ? 1'b0 : n638;
/* FF  8 11  1 */ assign n428 = n639;
/* FF  6 10  3 */ always @(posedge clk) if (1'b1) n259 <= 1'b0 ? 1'b0 : n640;
/* FF 11  9  4 */ always @(posedge clk) if (1'b1) n525 <= 1'b0 ? 1'b0 : n641;
/* FF  8 10  5 */ assign n425 = n642;
/* FF  5  4  0 */ always @(posedge clk) if (1'b1) n141 <= 1'b0 ? 1'b0 : n643;
/* FF  7  4  2 */ always @(posedge clk) if (1'b1) n301 <= 1'b0 ? 1'b0 : n644;
/* FF  9 11  3 */ assign n510 = n645;
/* FF  7  3  6 */ always @(posedge clk) if (1'b1) n299 <= 1'b0 ? 1'b0 : n646;
/* FF  4 10  3 */ always @(posedge clk) if (n2) n110 <= 1'b0 ? 1'b0 : n647;
/* FF  6  3  0 */ assign n65 = n648;
/* FF  6 14  0 */ assign n284 = n649;
/* FF  8 14  2 */ assign n452 = n650;
/* FF  8  3  2 */ always @(posedge clk) if (1'b1) n379 <= 1'b0 ? 1'b0 : n651;
/* FF  6  6  5 */ always @(posedge clk) if (1'b1) n232 <= 1'b0 ? 1'b0 : n652;
/* FF 11 12  5 */ assign n3 = n653;
/* FF  9  4  0 */ always @(posedge clk) if (1'b1) n461 <= 1'b0 ? 1'b0 : n654;
/* FF  5  7  1 */ always @(posedge clk) if (1'b1) n17 <= 1'b0 ? 1'b0 : n655;
/* FF  7 15  7 */ assign n375 = n656;
/* FF  4 11  4 */ always @(posedge clk) if (1'b1) n61 <= 1'b0 ? 1'b0 : n657;
/* FF  6 15  1 */ assign n208 = n658;
/* FF  7  7  3 */ always @(posedge clk) if (1'b1) n325 <= 1'b0 ? 1'b0 : n659;
/* FF  4  3  0 */ always @(posedge clk) if (1'b1) n79 <= 1'b0 ? 1'b0 : n660;
/* FF  9  7  5 */ always @(posedge clk) if (1'b1) n481 <= 1'b0 ? 1'b0 : n661;
/* FF  4 14  0 */ assign n662 = n663;
/* FF 11 13  6 */ always @(posedge clk) if (1'b1) n455 <= n3 ? 1'b0 : n665;
/* FF 12 12  0 */ always @(posedge clk) if (n532) d_vld <= 1'b0 ? 1'b0 : n666;
/* FF  5  8  2 */ always @(posedge clk) if (1'b1) n172 <= 1'b0 ? 1'b0 : n667;
/* FF  4 15  1 */ assign n39 = n668;
/* FF  4  4  1 */ always @(posedge clk) if (1'b1) n66 <= n4 ? 1'b0 : n669;
/* FF  7 11  0 */ assign n342 = n670;
/* FF  4  7  6 */ always @(posedge clk) if (1'b1) n92 <= 1'b0 ? 1'b0 : n671;
/* FF 11  6  3 */ always @(posedge clk) if (1'b1) n516 <= 1'b0 ? 1'b0 : n672;
/* FF  8 10  0 */ assign n420 = n673;
/* FF  6 10  7 */ always @(posedge clk) if (1'b1) n263 <= 1'b0 ? 1'b0 : n674;
/* FF  6 13  3 */ assign n278 = n675;
/* FF  7  3  1 */ always @(posedge clk) if (1'b1) n295 <= 1'b0 ? 1'b0 : n676;
/* FF  9 11  7 */ assign n336 = n677;
/* FF  9  3  3 */ always @(posedge clk) if (1'b1) n457 <= 1'b0 ? 1'b0 : n678;
/* FF  5  6  4 */ always @(posedge clk) if (1'b1) n14 <= 1'b0 ? 1'b0 : n679;
/* FF  6  3  4 */ always @(posedge clk) if (1'b1) n214 <= 1'b0 ? 1'b0 : n680;
/* FF  6 14  4 */ assign n286 = n681;
/* FF  8  3  6 */ always @(posedge clk) if (1'b1) n382 <= 1'b0 ? 1'b0 : n682;
/* FF  8 14  6 */ assign n454 = n683;
/* FF  5 15  0 */ always @(posedge clk) if (1'b1) n58 <= 1'b0 ? 1'b0 : n684;
/* FF  7 15  2 */ assign n373 = n685;
/* FF  9  4  4 */ always @(posedge clk) if (1'b1) n463 <= 1'b0 ? 1'b0 : n686;
/* FF  5  7  5 */ always @(posedge clk) if (1'b1) n163 <= 1'b0 ? 1'b0 : n687;
/* FF  9  7  0 */ assign n478 = n688;
/* FF  7  7  7 */ always @(posedge clk) if (1'b1) n329 <= 1'b0 ? 1'b0 : n689;
/* FF  4  3  4 */ always @(posedge clk) if (1'b1) n81 <= 1'b0 ? 1'b0 : n690;
/* FF  4 14  4 */ always @(posedge clk) if (n121) n126 <= rst ? 1'b0 : n691;
/* FF 11 13  1 */ assign n692 = n693;
/* FF 11  5  6 */ always @(posedge clk) if (1'b1) n29 <= 1'b0 ? 1'b0 : n694;
/* FF  6  9  1 */ always @(posedge clk) if (1'b1) n250 <= 1'b0 ? 1'b0 : n695;
/* FF  8  6  7 */ always @(posedge clk) if (1'b1) n401 <= 1'b0 ? 1'b0 : n696;
/* FF  7 14  6 */ assign n369 = n697;
/* FF  8 10  4 */ assign n424 = n698;
/* FF  6 13  7 */ assign n282 = n699;
/* FF  6  2  7 */ always @(posedge clk) if (1'b1) n210 <= n1 ? 1'b1 : n700;
/* FF  9 11  2 */ assign n509 = n701;
/* FF  5  3  3 */ always @(posedge clk) if (1'b1) n137 <= 1'b0 ? 1'b0 : n702;
/* FF  4 10  2 */ always @(posedge clk) if (n2) n109 <= 1'b0 ? 1'b0 : n703;
/* FF  8  3  1 */ assign n378 = n704;
/* FF  8 14  1 */ assign n451 = n705;
/* FF  6  6  4 */ always @(posedge clk) if (1'b1) n231 <= 1'b0 ? 1'b0 : n706;
/* FF 11 12  4 */ assign n533 = n707;
/* FF  5  7  0 */ assign n103 = n708;
/* FF  7 15  6 */ assign n374 = n709;
/* FF  7  7  2 */ always @(posedge clk) if (1'b1) n324 <= 1'b0 ? 1'b0 : n710;
/* FF  9  7  4 */ always @(posedge clk) if (1'b1) n332 <= 1'b0 ? 1'b0 : n711;
/* FF  5 10  2 */ always @(posedge clk) if (1'b1) n169 <= 1'b0 ? 1'b0 : n712;
/* FF  7 10  4 */ assign n340 = n713;
/* FF  8  6  2 */ assign n397 = n714;
/* FF  9 10  6 */ assign n501 = n715;
/* FF  6  9  5 */ always @(posedge clk) if (1'b1) n252 <= 1'b0 ? 1'b0 : n716;
/* FF  8  9  7 */ assign n209 = n717;
/* FF  7 14  1 */ assign n365 = n718;
/* FF 12  7  6 */ always @(posedge clk) if (1'b1) n536 <= 1'b0 ? 1'b0 : n719;
/* FF  6 10  6 */ always @(posedge clk) if (1'b1) n262 <= 1'b0 ? 1'b0 : n720;
/* FF  6 13  2 */ assign n277 = n721;
/* FF  9 11  6 */ assign n511 = n722;
/* FF  7  3  0 */ always @(posedge clk) if (1'b1) n294 <= 1'b0 ? 1'b0 : n723;
/* FF  5  3  7 */ always @(posedge clk) if (1'b1) n140 <= 1'b0 ? 1'b0 : n724;
/* FF  5  6  3 */ always @(posedge clk) if (1'b1) n155 <= 1'b0 ? 1'b0 : n725;
/* FF  4 10  6 */ always @(posedge clk) if (n2) n111 <= 1'b0 ? 1'b0 : n726;
/* FF  8 13  0 */ assign n442 = n727;
/* FF  6  5  3 */ always @(posedge clk) if (1'b1) n224 <= 1'b0 ? 1'b0 : n728;
/* FF  8  5  5 */ always @(posedge clk) if (1'b1) n393 <= 1'b0 ? 1'b0 : n729;
/* FF  5 10  6 */ always @(posedge clk) if (1'b1) n183 <= 1'b0 ? 1'b0 : n730;
/* FF  9 10  1 */ assign n503 = n731;
/* FF  6  9  0 */ always @(posedge clk) if (1'b1) n249 <= 1'b0 ? 1'b0 : n732;
/* FF  8  6  6 */ always @(posedge clk) if (1'b1) n400 <= 1'b0 ? 1'b0 : n733;
/* FF 11  7  5 */ always @(posedge clk) if (1'b1) n494 <= 1'b0 ? 1'b0 : n734;
/* FF 12  7  1 */ always @(posedge clk) if (1'b1) n535 <= 1'b0 ? 1'b0 : n735;
/* FF  6 10  1 */ always @(posedge clk) if (1'b1) n258 <= 1'b0 ? 1'b0 : n736;
/* FF  7 14  5 */ assign n368 = n737;
/* FF  8 10  3 */ assign n423 = n738;
/* FF  6 13  6 */ assign n281 = n739;
/* FF  9 11  1 */ assign n201 = n740;
/* FF  5  3  2 */ always @(posedge clk) if (1'b1) n136 <= 1'b0 ? 1'b0 : n741;
/* FF  7  3  4 */ always @(posedge clk) if (1'b1) n298 <= 1'b0 ? 1'b0 : n742;
/* FF  9  3  6 */ always @(posedge clk) if (1'b1) n460 <= 1'b0 ? 1'b0 : n743;
/* FF  5  6  7 */ always @(posedge clk) if (1'b1) n158 <= 1'b0 ? 1'b0 : n744;
/* FF  7  6  6 */ always @(posedge clk) if (1'b1) n319 <= 1'b0 ? 1'b0 : n745;
/* FF 11 12  3 */ assign n532 = n746;
/* FF  8 13  4 */ assign n83 = n747;
/* FF  8  5  0 */ always @(posedge clk) if (1'b1) n388 <= 1'b0 ? 1'b0 : n748;
/* FF  6  5  7 */ always @(posedge clk) if (1'b1) n228 <= 1'b0 ? 1'b0 : n749;
/* FF 11 11  7 */ always @(posedge clk) if (1'b1) n107 <= n123 ? 1'b1 : n750;
/* FF  5 10  1 */ always @(posedge clk) if (1'b1) n185 <= 1'b0 ? 1'b0 : n751;
/* FF  7 10  3 */ assign n339 = n752;
/* FF  8  6  1 */ assign n396 = n753;
/* FF  9 10  5 */ assign n506 = n754;
/* FF  6  9  4 */ always @(posedge clk) if (1'b1) n251 <= 1'b0 ? 1'b0 : n755;
/* FF  4  9  5 */ always @(posedge clk) if (1'b1) n25 <= n1 ? 1'b1 : n756;
/* FF  8  9  6 */ assign n8 = n757;
/* FF 11  7  0 */ always @(posedge clk) if (1'b1) n486 <= 1'b0 ? 1'b0 : n758;
/* FF  7 14  0 */ assign n364 = n759;
/* FF 11  8  1 */ always @(posedge clk) if (1'b1) n256 <= n1 ? 1'b1 : n760;
/* FF  6 12  5 */ assign n122 = n761;
/* FF  8 12  7 */ assign n440 = n762;
/* FF  7  6  1 */ always @(posedge clk) if (1'b1) n316 <= 1'b0 ? 1'b0 : n763;
/* FF  9  6  3 */ always @(posedge clk) if (1'b1) n69 <= 1'b0 ? 1'b0 : n764;
/* FF  5  9  4 */ always @(posedge clk) if (1'b1) n179 <= 1'b0 ? 1'b0 : n765;
/* FF  4 13  7 */ assign n121 = n766;
/* FF  2  5  1 */ always @(posedge clk) if (1'b1) n43 <= 1'b0 ? 1'b0 : n767;
/* FF  7  9  6 */ assign n334 = n768;
/* FF  6  5  2 */ always @(posedge clk) if (1'b1) n223 <= 1'b0 ? 1'b0 : n769;
/* FF  8  5  4 */ always @(posedge clk) if (1'b1) n392 <= 1'b0 ? 1'b0 : n770;
/* FF  5 10  5 */ always @(posedge clk) if (1'b1) \d_out[4]  <= 1'b0 ? 1'b0 : n771;
/* FF  9 10  0 */ assign n502 = n772;
/* FF  7 10  7 */ assign n106 = n773;
/* FF  8  9  1 */ assign n416 = n774;
/* FF 11  7  4 */ always @(posedge clk) if (1'b1) n520 <= 1'b0 ? 1'b0 : n775;
/* FF  4  6  3 */ always @(posedge clk) if (1'b1) n87 <= n4 ? 1'b0 : n776;
/* FF  5  5  2 */ always @(posedge clk) if (1'b1) n149 <= 1'b0 ? 1'b0 : n777;
/* FF  6 12  0 */ assign n271 = n778;
/* FF  7  5  4 */ always @(posedge clk) if (1'b1) n309 <= 1'b0 ? 1'b0 : n779;
/* FF  4 12  1 */ assign n116 = n780;
/* FF  8 12  2 */ assign n435 = n781;
/* FF  9  5  6 */ always @(posedge clk) if (1'b1) n471 <= 1'b0 ? 1'b0 : n782;
/* FF  8  4  7 */ always @(posedge clk) if (1'b1) n384 <= 1'b0 ? 1'b0 : n783;
/* FF  7  6  5 */ always @(posedge clk) if (1'b1) n241 <= 1'b0 ? 1'b0 : n784;
/* FF  8 13  3 */ assign n445 = n785;
/* FF  7  9  1 */ assign n168 = n786;
/* FF  9  6  7 */ always @(posedge clk) if (1'b1) n477 <= 1'b0 ? 1'b0 : n787;
/* FF  6  5  6 */ always @(posedge clk) if (1'b1) n227 <= 1'b0 ? 1'b0 : n788;
/* FF  5 10  0 */ always @(posedge clk) if (1'b1) n184 <= 1'b0 ? 1'b0 : n789;
/* FF  7 10  2 */ assign n338 = n790;
/* FF  9 10  4 */ assign n505 = n791;
/* FF  8  8  0 */ assign n406 = n792;
/* FF  2  8  6 */ always @(posedge clk) if (1'b1) n49 <= n1 ? 1'b1 : n793;
/* FF  6  8  7 */ always @(posedge clk) if (1'b1) n247 <= 1'b0 ? 1'b0 : n794;
/* FF  7 13  3 */ assign n358 = n795;
/* FF  9 13  5 */ always @(posedge clk) if (1'b1) n34 <= n3 ? 1'b0 : n796;
/* FF  5  5  6 */ always @(posedge clk) if (1'b1) n152 <= 1'b0 ? 1'b0 : n797;
/* FF  9  5  1 */ always @(posedge clk) if (1'b1) n466 <= 1'b0 ? 1'b0 : n798;
/* FF  6 12  4 */ assign n77 = n799;
/* FF  4 12  5 */ assign n75 = n800;
/* FF  6  4  0 */ always @(posedge clk) if (1'b1) n217 <= 1'b0 ? 1'b0 : n801;
/* FF  8 12  6 */ assign n439 = n802;
/* FF  8  4  2 */ always @(posedge clk) if (1'b1) n376 <= 1'b0 ? 1'b0 : n803;
/* FF  7  6  0 */ always @(posedge clk) if (1'b1) n315 <= 1'b0 ? 1'b0 : n804;
/* FF  9  6  2 */ always @(posedge clk) if (1'b1) n473 <= 1'b0 ? 1'b0 : n805;
/* FF  5  9  3 */ always @(posedge clk) if (1'b1) n178 <= 1'b0 ? 1'b0 : n806;
/* FF  7  9  5 */ assign n264 = n807;
/* FF  6  5  1 */ always @(posedge clk) if (1'b1) n222 <= 1'b0 ? 1'b0 : n808;
/* FF  8  5  3 */ always @(posedge clk) if (1'b1) n391 <= 1'b0 ? 1'b0 : n809;
/* FF  5 12  4 */ assign n199 = n810;
/* FF  7  1  6 */ assign n1 = n811;
/* FF  6  8  2 */ always @(posedge clk) if (1'b1) n20 <= 1'b0 ? 1'b0 : n812;
/* FF  7 12  6 */ assign n321 = n813;
/* FF  4  8  3 */ always @(posedge clk) if (1'b1) n97 <= 1'b0 ? 1'b0 : n814;
/* FF  8  8  4 */ always @(posedge clk) if (1'b1) \d_out[2]  <= 1'b0 ? 1'b0 : n815;
/* FF  2 11  6 */ always @(posedge clk) if (1'b1) n28 <= 1'b0 ? 1'b0 : n816;
/* FF  9 13  0 */ assign n512 = n817;
/* FF  5  5  1 */ always @(posedge clk) if (1'b1) n148 <= 1'b0 ? 1'b0 : n818;
/* FF  7 13  7 */ assign n195 = n819;
/* FF  8 12  1 */ assign n434 = n820;
/* FF  2 12  7 */ always @(posedge clk) if (1'b1) n57 <= 1'b0 ? 1'b0 : n821;
/* FF  9  5  5 */ always @(posedge clk) if (1'b1) n470 <= 1'b0 ? 1'b0 : n822;
/* FF  6  4  4 */ always @(posedge clk) if (1'b1) n219 <= 1'b0 ? 1'b0 : n823;
/* FF  6  7  6 */ always @(posedge clk) if (1'b1) n239 <= 1'b0 ? 1'b0 : n824;
/* FF  9  6  6 */ always @(posedge clk) if (1'b1) n476 <= 1'b0 ? 1'b0 : n825;
/* FF  7  9  0 */ assign n167 = n826;
/* FF 11 11  5 */ always @(posedge clk) if (1'b1) n42 <= n123 ? 1'b0 : n827;
/* FF 11  3  1 */ always @(posedge clk) if (1'b1) \d_out[1]  <= 1'b0 ? 1'b0 : n828;
/* FF  6 11  3 */ assign n268 = n829;
/* FF  8 11  5 */ assign n275 = n830;
/* FF  7 12  1 */ assign n283 = n831;
/* FF  2  8  5 */ assign n48 = n832;
/* FF  5  4  4 */ always @(posedge clk) if (1'b1) \d_out[5]  <= 1'b0 ? 1'b0 : n833;
/* FF  6  8  6 */ always @(posedge clk) if (1'b1) n246 <= 1'b0 ? 1'b0 : n834;
/* FF  4  8  7 */ always @(posedge clk) if (1'b1) n100 <= 1'b0 ? 1'b0 : n835;
/* FF  7  4  6 */ always @(posedge clk) if (1'b1) n305 <= 1'b0 ? 1'b0 : n836;
/* FF  7 13  2 */ assign n357 = n837;
/* FF  5  5  5 */ always @(posedge clk) if (1'b1) n151 <= 1'b0 ? 1'b0 : n838;
/* FF  9  5  0 */ always @(posedge clk) if (1'b1) n465 <= 1'b0 ? 1'b0 : n839;
/* FF  2 12  2 */ always @(posedge clk) if (1'b1) n32 <= 1'b0 ? 1'b0 : n840;
/* FF  7  5  7 */ always @(posedge clk) if (1'b1) n312 <= 1'b0 ? 1'b0 : n841;
/* FF  4 12  4 */ assign n74 = n842;
/* FF  6  7  1 */ assign n235 = n843;
/* FF  8  7  3 */ always @(posedge clk) if (1'b1) n50 <= 1'b0 ? 1'b0 : n844;
/* FF  5  8  6 */ always @(posedge clk) if (1'b1) n175 <= 1'b0 ? 1'b0 : n845;
/* FF  9  8  1 */ always @(posedge clk) if (1'b1) n488 <= 1'b0 ? 1'b0 : n846;
/* FF  4 15  5 */ assign n64 = n847;
/* FF  7 11  4 */ assign n346 = n848;
/* FF  4  7  1 */ always @(posedge clk) if (1'b1) n90 <= 1'b0 ? 1'b0 : n849;
/* FF  8 11  0 */ assign n418 = n850;
/* FF  6 11  7 */ always @(posedge clk) if (n2) n270 <= 1'b0 ? 1'b0 : n851;
/* FF 11  6  7 */ always @(posedge clk) if (1'b1) n484 <= 1'b0 ? 1'b0 : n852;
/* FF 11  9  3 */ always @(posedge clk) if (1'b1) n187 <= 1'b0 ? 1'b0 : n853;
/* FF  5 12  3 */ assign n198 = n854;
/* FF  7 12  5 */ assign n204 = n855;
/* FF  6  8  1 */ always @(posedge clk) if (1'b1) n245 <= 1'b0 ? 1'b0 : n856;
/* FF  4  8  2 */ always @(posedge clk) if (1'b1) n96 <= 1'b0 ? 1'b0 : n857;
/* FF  7  4  1 */ assign n300 = n858;
/* FF  8  8  3 */ always @(posedge clk) if (1'b1) n410 <= 1'b0 ? 1'b0 : n859;
/* FF 11 10  4 */ always @(posedge clk) if (1'b1) n15 <= 1'b0 ? 1'b0 : n860;
/* FF  5  5  0 */ always @(posedge clk) if (1'b1) n147 <= 1'b0 ? 1'b0 : n861;
/* FF  7  5  2 */ always @(posedge clk) if (1'b1) n308 <= 1'b0 ? 1'b0 : n862;
/* FF  9  5  4 */ always @(posedge clk) if (1'b1) n469 <= 1'b0 ? 1'b0 : n863;
/* FF  2  4  2 */ always @(posedge clk) if (1'b1) n11 <= 1'b0 ? 1'b0 : n864;
/* FF  4 11  3 */ always @(posedge clk) if (1'b1) n108 <= 1'b0 ? 1'b0 : n865;
/* FF  6 15  0 */ assign n289 = n866;
/* FF  6  7  5 */ always @(posedge clk) if (1'b1) n238 <= 1'b0 ? 1'b0 : n867;
/* FF  8  7  7 */ always @(posedge clk) if (1'b1) n405 <= 1'b0 ? 1'b0 : n868;
/* FF 11 13  5 */ always @(posedge clk) if (1'b1) n188 <= n3 ? 1'b0 : n869;
/* FF  5  8  1 */ always @(posedge clk) if (1'b1) n171 <= 1'b0 ? 1'b0 : n870;
/* FF  4 15  0 */ assign n128 = n871;
/* FF  9  8  5 */ always @(posedge clk) if (1'b1) n491 <= 1'b0 ? 1'b0 : n872;
/* FF  5 11  6 */ always @(posedge clk) if (1'b1) n194 <= n4 ? 1'b0 : n873;
/* FF  2  7  3 */ always @(posedge clk) if (1'b1) n18 <= 1'b0 ? 1'b0 : n874;
/* FF  4  7  5 */ always @(posedge clk) if (1'b1) n51 <= 1'b0 ? 1'b0 : n875;
/* FF  6 11  2 */ assign n267 = n876;
/* FF  8 11  4 */ assign n430 = n877;
/* FF 11  9  7 */ always @(posedge clk) if (1'b1) n528 <= 1'b0 ? 1'b0 : n878;
/* FF  7 12  0 */ assign n349 = n879;
/* FF  5  4  3 */ always @(posedge clk) if (1'b1) n143 <= 1'b0 ? 1'b0 : n880;
/* FF  4  8  6 */ always @(posedge clk) if (1'b1) n54 <= 1'b0 ? 1'b0 : n881;
/* FF  7  4  5 */ always @(posedge clk) if (1'b1) n304 <= 1'b0 ? 1'b0 : n882;
/* FF  6  3  3 */ always @(posedge clk) if (1'b1) n213 <= 1'b0 ? 1'b0 : n883;
/* FF  8 14  5 */ assign n441 = n884;
/* FF  7 15  1 */ assign n372 = n885;
/* FF  5  7  4 */ always @(posedge clk) if (1'b1) n162 <= 1'b0 ? 1'b0 : n886;
/* FF  6 15  4 */ assign n4 = n887;
/* FF  7  7  6 */ always @(posedge clk) if (1'b1) n328 <= 1'b0 ? 1'b0 : n888;
/* FF  4  3  3 */ always @(posedge clk) if (1'b1) n80 <= 1'b0 ? 1'b0 : n889;
/* FF  6  7  0 */ assign n234 = n890;
/* FF  4 14  3 */ always @(posedge clk) if (n121) n125 <= rst ? 1'b0 : n891;
/* FF  8  7  2 */ always @(posedge clk) if (1'b1) n72 <= 1'b0 ? 1'b0 : n892;
/* FF 11 13  0 */ assign n893 = n894;
/* FF 11  5  5 */ always @(posedge clk) if (1'b1) n515 <= 1'b0 ? 1'b0 : n896;
/* FF  5  8  5 */ always @(posedge clk) if (1'b1) n70 <= 1'b0 ? 1'b0 : n897;
/* FF  9  8  0 */ always @(posedge clk) if (1'b1) n487 <= 1'b0 ? 1'b0 : n898;
/* FF  2 15  2 */ always @(posedge clk) if (1'b1) n52 <= 1'b0 ? 1'b0 : n899;
/* FF  5 11  1 */ assign n191 = n900;
/* FF  4 15  4 */ assign n63 = n901;
/* FF  7 11  3 */ assign n345 = n902;
/* FF  4  7  0 */ always @(posedge clk) if (1'b1) n89 <= 1'b0 ? 1'b0 : n903;
/* FF  2  7  7 */ always @(posedge clk) if (1'b1) n46 <= 1'b0 ? 1'b0 : n904;
/* FF 11  6  6 */ always @(posedge clk) if (1'b1) n518 <= 1'b0 ? 1'b0 : n905;
/* FF 11  9  2 */ always @(posedge clk) if (1'b1) n524 <= 1'b0 ? 1'b0 : n906;
/* FF  7 12  4 */ assign n350 = n907;
/* FF  4  8  1 */ always @(posedge clk) if (1'b1) n95 <= 1'b0 ? 1'b0 : n908;
/* FF  7  4  0 */ assign n159 = n909;
/* FF  8 14  0 */ assign n449 = n910;
/* FF  8  3  0 */ assign n377 = n911;
/* FF  6  3  7 */ always @(posedge clk) if (1'b1) n216 <= 1'b0 ? 1'b0 : n912;
/* FF  6 14  7 */ assign n132 = n913;
/* FF  4 11  2 */ assign n114 = n914;
/* FF  7  7  1 */ assign n323 = n915;
/* FF  9  4  7 */ always @(posedge clk) if (1'b1) n313 <= 1'b0 ? 1'b0 : n916;
/* FF  9  7  3 */ always @(posedge clk) if (1'b1) n73 <= 1'b0 ? 1'b0 : n917;
/* FF  4  3  7 */ always @(posedge clk) if (1'b1) n82 <= 1'b0 ? 1'b0 : n918;
/* FF  6  7  4 */ always @(posedge clk) if (1'b1) n237 <= 1'b0 ? 1'b0 : n919;
/* FF  8  7  6 */ always @(posedge clk) if (1'b1) n404 <= 1'b0 ? 1'b0 : n920;
/* FF 11 13  4 */ always @(posedge clk) if (1'b1) n433 <= n3 ? 1'b0 : n921;
/* FF 11  5  0 */ assign n101 = n922;
/* FF  5  8  0 */ always @(posedge clk) if (1'b1) n170 <= 1'b0 ? 1'b0 : n923;
/* FF  9  8  4 */ always @(posedge clk) if (1'b1) n490 <= 1'b0 ? 1'b0 : n924;
/* FF  2 15  6 */ always @(posedge clk) if (1'b1) n38 <= 1'b0 ? 1'b0 : n925;
/* FF  2  7  2 */ always @(posedge clk) if (1'b1) n19 <= 1'b0 ? 1'b0 : n926;
/* FF 11  6  1 */ always @(posedge clk) if (1'b1) n104 <= 1'b0 ? 1'b0 : n927;
/* FF  5 14  7 */ assign n189 = n928;
/* FF  6 10  5 */ always @(posedge clk) if (1'b1) n261 <= 1'b0 ? 1'b0 : n929;
/* FF 11  9  6 */ always @(posedge clk) if (1'b1) n527 <= 1'b0 ? 1'b0 : n930;
/* FF  8 10  7 */ assign n426 = n931;
/* FF  9 11  5 */ assign n353 = n932;
/* FF  5  3  6 */ always @(posedge clk) if (1'b1) n139 <= 1'b0 ? 1'b0 : n933;
/* FF  4 10  5 */ always @(posedge clk) if (n2) n60 <= 1'b0 ? 1'b0 : n934;
/* FF  6 14  2 */ assign n36 = n935;
/* FF  6  3  2 */ always @(posedge clk) if (1'b1) n212 <= 1'b0 ? 1'b0 : n936;
/* FF  8 14  4 */ assign n450 = n937;
/* FF  8  3  4 */ always @(posedge clk) if (1'b1) n381 <= 1'b0 ? 1'b0 : n938;
/* FF  7 15  0 */ assign n362 = n939;
/* FF 11  4  3 */ always @(posedge clk) if (1'b1) n514 <= n4 ? 1'b0 : n940;
/* FF  5 15  7 */ always @(posedge clk) if (1'b1) n205 <= 1'b0 ? 1'b0 : n941;
/* FF  5  7  3 */ always @(posedge clk) if (1'b1) n161 <= 1'b0 ? 1'b0 : n942;
/* FF  4 11  6 */ always @(posedge clk) if (1'b1) n115 <= 1'b0 ? 1'b0 : n943;
/* FF  7  7  5 */ always @(posedge clk) if (1'b1) n327 <= 1'b0 ? 1'b0 : n944;
/* FF  4  3  2 */ always @(posedge clk) if (1'b1) n12 <= 1'b0 ? 1'b0 : n945;
/* FF  4 14  2 */ always @(posedge clk) if (n121) n124 <= rst ? 1'b0 : n946;
/* FF  9  7  7 */ always @(posedge clk) if (1'b1) n483 <= 1'b0 ? 1'b0 : n947;
/* FF  8  7  1 */ always @(posedge clk) if (1'b1) n403 <= 1'b0 ? 1'b0 : n948;
/* FF  8  6  5 */ always @(posedge clk) if (1'b1) \d_out[0]  <= 1'b0 ? 1'b0 : n949;
/* FF  5 11  0 */ assign n190 = n950;
/* FF  7 11  2 */ assign n344 = n951;
/* FF  7 14  4 */ assign n367 = n952;
/* FF  6 10  0 */ always @(posedge clk) if (1'b1) n257 <= 1'b0 ? 1'b0 : n953;
/* FF 11  9  1 */ always @(posedge clk) if (1'b1) n523 <= 1'b0 ? 1'b0 : n954;
/* FF  8 10  2 */ assign n422 = n955;
/* FF  6 13  5 */ assign n280 = n956;
/* FF  9 11  0 */ assign n508 = n957;
/* FF  5  3  1 */ always @(posedge clk) if (1'b1) n135 <= 1'b0 ? 1'b0 : n958;
/* FF  7  3  3 */ always @(posedge clk) if (1'b1) n297 <= 1'b0 ? 1'b0 : n959;
/* FF  9  3  5 */ always @(posedge clk) if (1'b1) n459 <= 1'b0 ? 1'b0 : n960;
/* FF  5  6  6 */ always @(posedge clk) if (1'b1) n157 <= 1'b0 ? 1'b0 : n961;
/* FF  6 14  6 */ assign n288 = n962;
/* FF  6  6  2 */ always @(posedge clk) if (1'b1) n230 <= 1'b0 ? 1'b0 : n963;
/* FF  5 15  2 */ always @(posedge clk) if (1'b1) n2 <= 1'b0 ? 1'b0 : n964;
/* FF  7 15  4 */ assign n363 = n965;
/* FF  7  7  0 */ assign n322 = n966;
/* FF  9  4  6 */ always @(posedge clk) if (1'b1) n464 <= 1'b0 ? 1'b0 : n967;
/* FF  5  7  7 */ always @(posedge clk) if (1'b1) n102 <= 1'b0 ? 1'b0 : n968;
/* FF  9  7  2 */ assign n480 = n969;
/* FF 11 13  3 */ always @(posedge clk) if (1'b1) n534 <= n3 ? 1'b0 : n970;
/* FF  6  9  3 */ always @(posedge clk) if (1'b1) n243 <= 1'b0 ? 1'b0 : n971;
/* FF  8  9  5 */ assign n407 = n972;
/* FF  9 14  1 */ always @(posedge clk) if (1'b1) n123 <= 1'b0 ? 1'b0 : n973;
/* FF  4  6  7 */ always @(posedge clk) if (1'b1) n85 <= n4 ? 1'b0 : n974;
/* FF  6 10  4 */ always @(posedge clk) if (1'b1) n260 <= 1'b0 ? 1'b0 : n975;
/* FF  6 13  0 */ assign n276 = n976;
/* FF  8 10  6 */ assign n419 = n977;
/* FF  9 11  4 */ assign n352 = n978;
/* FF  5  3  5 */ always @(posedge clk) if (1'b1) n138 <= 1'b0 ? 1'b0 : n979;
/* FF  5  6  1 */ always @(posedge clk) if (1'b1) n154 <= 1'b0 ? 1'b0 : n980;
/* FF  8 14  3 */ assign n453 = n981;
/* FF  8 13  7 */ assign n448 = n982;
/* FF  9  4  1 */ always @(posedge clk) if (1'b1) n462 <= 1'b0 ? 1'b0 : n983;
/* FF  5  7  2 */ always @(posedge clk) if (1'b1) n71 <= 1'b0 ? 1'b0 : n984;
/* FF  7  7  4 */ always @(posedge clk) if (1'b1) n326 <= 1'b0 ? 1'b0 : n985;
/* FF  4  3  1 */ always @(posedge clk) if (1'b1) \d_out[6]  <= 1'b0 ? 1'b0 : n986;
/* FF  4 14  1 */ assign n987 = n988;
/* FF  9  7  6 */ always @(posedge clk) if (1'b1) n482 <= 1'b0 ? 1'b0 : n989;
/* FF  5 10  4 */ always @(posedge clk) if (1'b1) n176 <= 1'b0 ? 1'b0 : n990;
/* FF  7 10  6 */ assign n10 = n991;
/* FF  8  6  4 */ always @(posedge clk) if (1'b1) n398 <= 1'b0 ? 1'b0 : n992;
/* FF  8  9  0 */ assign n415 = n993;
/* FF  6  9  7 */ always @(posedge clk) if (1'b1) n254 <= 1'b0 ? 1'b0 : n994;
/* FF  7 14  3 */ assign n354 = n995;
/* FF  8 10  1 */ assign n421 = n996;
/* FF  6 13  4 */ assign n279 = n997;
/* FF  7  3  2 */ always @(posedge clk) if (1'b1) n296 <= 1'b0 ? 1'b0 : n998;
/* FF  9  3  4 */ always @(posedge clk) if (1'b1) n458 <= 1'b0 ? 1'b0 : n999;
/* FF  2 10  6 */ always @(posedge clk) if (1'b1) n26 <= 1'b0 ? 1'b0 : n1000;
/* FF  5  6  5 */ always @(posedge clk) if (1'b1) n156 <= 1'b0 ? 1'b0 : n1001;
/* FF  7  6  4 */ always @(posedge clk) if (1'b1) n318 <= 1'b0 ? 1'b0 : n1002;
/* FF 11 12  1 */ assign n531 = n1003;
/* FF  8 13  2 */ assign n444 = n1004;
/* FF  5  9  7 */ always @(posedge clk) if (1'b1) n182 <= 1'b0 ? 1'b0 : n1005;
/* FF  1 12  0 */ always @(posedge clk) if (1'b1) n27 <= n4 ? 1'b0 : n1006;
/* FF  6  5  5 */ always @(posedge clk) if (1'b1) n226 <= 1'b0 ? 1'b0 : n1007;
/* FF  8  5  7 */ always @(posedge clk) if (1'b1) n395 <= 1'b0 ? 1'b0 : n1008;
/* FF  7 10  1 */ assign n337 = n1009;
/* FF  9 10  3 */ assign n348 = n1010;
/* FF  6  9  2 */ always @(posedge clk) if (1'b1) n24 <= 1'b0 ? 1'b0 : n1011;
/* FF  8  9  4 */ assign n417 = n1012;
/* FF 11  7  7 */ always @(posedge clk) if (1'b1) n521 <= 1'b0 ? 1'b0 : n1013;
/* FF  2  6  4 */ always @(posedge clk) if (1'b1) n13 <= n1 ? 1'b1 : n1014;
/* FF 12  7  3 */ always @(posedge clk) if (1'b1) n248 <= 1'b0 ? 1'b0 : n1015;
/* FF  7 14  7 */ assign n370 = n1016;
/* FF  6 12  3 */ assign n6 = n1017;
/* FF  8 12  5 */ assign n438 = n1018;
/* FF  5  6  0 */ assign n47 = n1019;
/* FF  9  6  1 */ always @(posedge clk) if (1'b1) n165 <= 1'b0 ? 1'b0 : n1020;
/* FF  5  9  2 */ always @(posedge clk) if (1'b1) n177 <= 1'b0 ? 1'b0 : n1021;
/* FF  7  9  4 */ assign n333 = n1022;
/* FF  6  5  0 */ always @(posedge clk) if (1'b1) n221 <= 1'b0 ? 1'b0 : n1023;
/* FF  8 13  6 */ assign n447 = n1024;
/* FF 11 11  0 */ assign n529 = n1025;
/* FF  9  9  6 */ always @(posedge clk) if (1'b1) n500 <= 1'b0 ? 1'b0 : n1026;
/* FF  8  5  2 */ always @(posedge clk) if (1'b1) n390 <= 1'b0 ? 1'b0 : n1027;
/* FF  7 10  5 */ assign n341 = n1028;
/* FF  9 10  7 */ assign n507 = n1029;
/* FF  6  9  6 */ always @(posedge clk) if (1'b1) n253 <= 1'b0 ? 1'b0 : n1030;
/* FF  4  9  7 */ always @(posedge clk) if (1'b1) n105 <= n1 ? 1'b1 : n1031;
/* FF 11  7  2 */ always @(posedge clk) if (1'b1) n519 <= 1'b0 ? 1'b0 : n1032;
/* FF  4  6  1 */ always @(posedge clk) if (1'b1) n86 <= n4 ? 1'b1 : n1033;
/* FF  7 14  2 */ assign n366 = n1034;
/* FF  7 13  6 */ assign n361 = n1035;
/* FF 11  8  3 */ always @(posedge clk) if (1'b1) n522 <= n1 ? 1'b1 : n1036;
/* FF  8 12  0 */ assign n88 = n1037;
/* FF  2 12  6 */ always @(posedge clk) if (1'b1) n56 <= 1'b0 ? 1'b0 : n1038;
/* FF  6 12  7 */ assign n274 = n1039;
/* FF  6  4  3 */ always @(posedge clk) if (1'b1) n160 <= 1'b0 ? 1'b0 : n1040;
/* FF  8  4  5 */ always @(posedge clk) if (1'b1) n387 <= 1'b0 ? 1'b0 : n1041;
/* FF  7  6  3 */ always @(posedge clk) if (1'b1) n317 <= 1'b0 ? 1'b0 : n1042;
/* FF  9  6  5 */ always @(posedge clk) if (1'b1) n475 <= 1'b0 ? 1'b0 : n1043;
/* FF  2 13  7 */ assign n35 = n1044;
/* FF  5  9  6 */ always @(posedge clk) if (1'b1) n181 <= 1'b0 ? 1'b0 : n1045;
/* FF  8 13  1 */ assign n443 = n1046;
/* FF  9  9  1 */ assign n497 = n1047;
/* FF  6  5  4 */ always @(posedge clk) if (1'b1) n225 <= 1'b0 ? 1'b0 : n1048;
/* FF  8  5  6 */ always @(posedge clk) if (1'b1) n394 <= 1'b0 ? 1'b0 : n1049;
/* FF 11 11  4 */ always @(posedge clk) if (1'b1) n7 <= n123 ? 1'b1 : n1050;
/* FF  9 10  2 */ assign n504 = n1051;
/* FF  8  9  3 */ assign n53 = n1052;
/* FF 11  7  6 */ always @(posedge clk) if (1'b1) n495 <= 1'b0 ? 1'b0 : n1053;
/* FF  8  8  7 */ always @(posedge clk) if (1'b1) n414 <= 1'b0 ? 1'b0 : n1054;
/* FF  7 13  1 */ assign n356 = n1055;
/* FF  9 13  3 */ always @(posedge clk) if (1'b1) n76 <= n3 ? 1'b0 : n1056;
/* FF  2 12  1 */ assign n31 = n1057;
/* FF  7  5  6 */ always @(posedge clk) if (1'b1) n311 <= 1'b0 ? 1'b0 : n1058;
/* FF  6 12  2 */ assign n273 = n1059;
/* FF  4 12  3 */ assign n118 = n1060;
/* FF  8 12  4 */ assign n437 = n1061;
/* FF  8  4  0 */ always @(posedge clk) if (1'b1) n385 <= 1'b0 ? 1'b0 : n1062;
/* FF  6  4  7 */ always @(posedge clk) if (1'b1) \d_out[3]  <= 1'b0 ? 1'b0 : n1063;
/* FF  9  6  0 */ assign n472 = n1064;
/* FF  5  9  1 */ assign n112 = n1065;
/* FF  7  6  7 */ always @(posedge clk) if (1'b1) n320 <= 1'b0 ? 1'b0 : n1066;
/* FF  7  9  3 */ assign n242 = n1067;
/* FF  8 13  5 */ assign n446 = n1068;
/* FF  9  9  5 */ assign n499 = n1069;
/* FF  8  5  1 */ always @(posedge clk) if (1'b1) n389 <= 1'b0 ? 1'b0 : n1070;
/* FF  6 11  6 */ assign n265 = n1071;
/* FF  6  8  0 */ always @(posedge clk) if (1'b1) n244 <= 1'b0 ? 1'b0 : n1072;
/* FF  8  8  2 */ always @(posedge clk) if (1'b1) n409 <= 1'b0 ? 1'b0 : n1073;
/* FF  5  4  7 */ always @(posedge clk) if (1'b1) n146 <= 1'b0 ? 1'b0 : n1074;
/* FF  7 13  5 */ assign n360 = n1075;
/* FF  7  5  1 */ assign n68 = n1076;
/* FF 12  9  6 */ always @(posedge clk) if (1'b1) n537 <= n1 ? 1'b1 : n1077;
/* FF  9  5  3 */ always @(posedge clk) if (1'b1) n468 <= 1'b0 ? 1'b0 : n1078;
/* FF  6 12  6 */ assign n133 = n1079;
/* FF  4 12  7 */ always @(posedge clk) if (n2) n120 <= 1'b0 ? 1'b0 : n1080;
/* FF  6  4  2 */ always @(posedge clk) if (1'b1) n218 <= 1'b0 ? 1'b0 : n1081;
/* FF  8  4  4 */ always @(posedge clk) if (1'b1) n386 <= 1'b0 ? 1'b0 : n1082;
/* FF  7  6  2 */ always @(posedge clk) if (1'b1) n314 <= 1'b0 ? 1'b0 : n1083;
/* FF  9  6  4 */ always @(posedge clk) if (1'b1) n474 <= 1'b0 ? 1'b0 : n1084;
/* FF  5  9  5 */ always @(posedge clk) if (1'b1) n180 <= 1'b0 ? 1'b0 : n1085;
/* FF  9  9  0 */ assign n496 = n1086;
/* FF  2  5  2 */ always @(posedge clk) if (1'b1) n44 <= 1'b0 ? 1'b0 : n1087;
/* FF  7  9  7 */ always @(posedge clk) if (1'b1) n335 <= n4 ? 1'b1 : n1088;
/* FF  6 11  1 */ assign n266 = n1089;
/* FF  8 11  3 */ assign n429 = n1090;

// Warning: unmatched port '\d_in[7] '
// Warning: unmatched port '\d_in[5] '
// Warning: unmatched port '\d_in[6] '
// Warning: unmatched port '\d_in[3] '
// Warning: unmatched port '\d_in[0] '
// Warning: unmatched port '\d_in[4] '
// Warning: unmatched port '\d_in[1] '
// Warning: unmatched port '\d_in[2] '

endmodule

