// Reading file 'aes_trojan.asc'..

module chip (input clk, output d_vld, input rst, output \d_out[6] , output \d_out[7] , output \d_out[5] , output \d_out[4] , output \d_out[3] , output \d_out[0] , output \d_out[2] , output \d_out[1] , input io_10_17_1);

wire n1;
// (0, 0, 'glb_netwk_0')
// (2, 3, 'lutff_global/s_r')
// (2, 4, 'lutff_global/s_r')
// (6, 2, 'neigh_op_tnr_2')
// (6, 3, 'neigh_op_rgt_2')
// (6, 4, 'neigh_op_bnr_2')
// (7, 0, 'fabout')
// (7, 0, 'local_g1_0')
// (7, 0, 'span12_vert_8')
// (7, 1, 'sp12_v_b_8')
// (7, 2, 'neigh_op_top_2')
// (7, 2, 'sp12_v_b_7')
// (7, 3, 'lutff_2/out')
// (7, 3, 'sp12_v_b_4')
// (7, 4, 'neigh_op_bot_2')
// (7, 4, 'sp12_v_b_3')
// (7, 5, 'sp12_v_b_0')
// (8, 2, 'neigh_op_tnl_2')
// (8, 3, 'neigh_op_lft_2')
// (8, 4, 'neigh_op_bnl_2')

wire n2;
// (0, 0, 'glb_netwk_2')
// (1, 10, 'lutff_global/s_r')
// (2, 6, 'lutff_global/s_r')
// (5, 5, 'lutff_global/s_r')
// (7, 4, 'lutff_global/s_r')
// (7, 6, 'lutff_global/s_r')
// (9, 3, 'glb2local_0')
// (9, 3, 'local_g0_4')
// (9, 3, 'lutff_5/in_3')
// (10, 7, 'neigh_op_tnr_1')
// (10, 8, 'neigh_op_rgt_1')
// (10, 8, 'sp4_h_r_7')
// (10, 9, 'neigh_op_bnr_1')
// (11, 7, 'neigh_op_top_1')
// (11, 8, 'lutff_1/out')
// (11, 8, 'lutff_global/s_r')
// (11, 8, 'sp4_h_r_18')
// (11, 9, 'neigh_op_bot_1')
// (12, 7, 'neigh_op_tnl_1')
// (12, 8, 'neigh_op_lft_1')
// (12, 8, 'sp4_h_r_31')
// (12, 9, 'neigh_op_bnl_1')
// (13, 8, 'span4_horz_31')
// (13, 8, 'span4_vert_t_13')
// (13, 9, 'fabout')
// (13, 9, 'local_g0_5')
// (13, 9, 'span4_vert_b_13')
// (13, 10, 'span4_vert_b_9')
// (13, 11, 'span4_vert_b_5')
// (13, 12, 'span4_vert_b_1')

wire clk;
// (0, 0, 'glb_netwk_3')
// (0, 5, 'span4_vert_t_14')
// (0, 6, 'span4_vert_b_14')
// (0, 7, 'span4_vert_b_10')
// (0, 8, 'io_1/D_IN_0')
// (0, 8, 'io_1/PAD')
// (0, 8, 'span4_vert_b_6')
// (0, 9, 'fabout')
// (0, 9, 'local_g1_2')
// (0, 9, 'span4_vert_b_2')
// (1, 7, 'neigh_op_tnl_2')
// (1, 7, 'neigh_op_tnl_6')
// (1, 8, 'lutff_global/clk')
// (1, 8, 'neigh_op_lft_2')
// (1, 8, 'neigh_op_lft_6')
// (1, 9, 'neigh_op_bnl_2')
// (1, 9, 'neigh_op_bnl_6')
// (1, 10, 'lutff_global/clk')
// (1, 12, 'lutff_global/clk')
// (2, 3, 'lutff_global/clk')
// (2, 4, 'lutff_global/clk')
// (2, 5, 'lutff_global/clk')
// (2, 6, 'lutff_global/clk')
// (2, 7, 'lutff_global/clk')
// (2, 8, 'lutff_global/clk')
// (2, 9, 'lutff_global/clk')
// (2, 10, 'lutff_global/clk')
// (2, 11, 'lutff_global/clk')
// (2, 12, 'lutff_global/clk')
// (2, 13, 'lutff_global/clk')
// (2, 14, 'lutff_global/clk')
// (4, 4, 'lutff_global/clk')
// (4, 5, 'lutff_global/clk')
// (4, 6, 'lutff_global/clk')
// (4, 7, 'lutff_global/clk')
// (4, 8, 'lutff_global/clk')
// (4, 9, 'lutff_global/clk')
// (4, 11, 'lutff_global/clk')
// (4, 12, 'lutff_global/clk')
// (4, 13, 'lutff_global/clk')
// (4, 14, 'lutff_global/clk')
// (5, 3, 'lutff_global/clk')
// (5, 4, 'lutff_global/clk')
// (5, 5, 'lutff_global/clk')
// (5, 7, 'lutff_global/clk')
// (5, 8, 'lutff_global/clk')
// (5, 9, 'lutff_global/clk')
// (5, 10, 'lutff_global/clk')
// (5, 11, 'lutff_global/clk')
// (5, 12, 'lutff_global/clk')
// (5, 13, 'lutff_global/clk')
// (5, 14, 'lutff_global/clk')
// (6, 7, 'lutff_global/clk')
// (6, 8, 'lutff_global/clk')
// (6, 9, 'lutff_global/clk')
// (6, 10, 'lutff_global/clk')
// (6, 11, 'lutff_global/clk')
// (6, 12, 'lutff_global/clk')
// (6, 13, 'lutff_global/clk')
// (6, 14, 'lutff_global/clk')
// (7, 4, 'lutff_global/clk')
// (7, 6, 'lutff_global/clk')
// (7, 7, 'lutff_global/clk')
// (7, 8, 'lutff_global/clk')
// (7, 9, 'lutff_global/clk')
// (7, 10, 'lutff_global/clk')
// (7, 11, 'lutff_global/clk')
// (7, 12, 'lutff_global/clk')
// (7, 13, 'lutff_global/clk')
// (7, 14, 'lutff_global/clk')
// (8, 5, 'lutff_global/clk')
// (8, 6, 'lutff_global/clk')
// (8, 7, 'lutff_global/clk')
// (8, 8, 'lutff_global/clk')
// (8, 9, 'lutff_global/clk')
// (8, 10, 'lutff_global/clk')
// (8, 11, 'lutff_global/clk')
// (8, 12, 'lutff_global/clk')
// (8, 13, 'lutff_global/clk')
// (8, 14, 'lutff_global/clk')
// (8, 15, 'lutff_global/clk')
// (9, 4, 'lutff_global/clk')
// (9, 5, 'lutff_global/clk')
// (9, 6, 'lutff_global/clk')
// (9, 7, 'lutff_global/clk')
// (9, 8, 'lutff_global/clk')
// (9, 9, 'lutff_global/clk')
// (9, 10, 'lutff_global/clk')
// (9, 11, 'lutff_global/clk')
// (9, 12, 'lutff_global/clk')
// (9, 13, 'lutff_global/clk')
// (11, 3, 'lutff_global/clk')
// (11, 4, 'lutff_global/clk')
// (11, 5, 'lutff_global/clk')
// (11, 6, 'lutff_global/clk')
// (11, 7, 'lutff_global/clk')
// (11, 8, 'lutff_global/clk')
// (11, 9, 'lutff_global/clk')
// (11, 11, 'lutff_global/clk')
// (11, 12, 'lutff_global/clk')
// (11, 13, 'lutff_global/clk')

wire n4;
// (0, 0, 'glb_netwk_6')
// (0, 7, 'logic_op_tnr_0')
// (0, 8, 'fabout')
// (0, 8, 'local_g1_0')
// (0, 8, 'logic_op_rgt_0')
// (0, 9, 'logic_op_bnr_0')
// (1, 7, 'neigh_op_top_0')
// (1, 8, 'lutff_0/out')
// (1, 8, 'lutff_global/s_r')
// (1, 9, 'neigh_op_bot_0')
// (2, 7, 'neigh_op_tnl_0')
// (2, 8, 'neigh_op_lft_0')
// (2, 9, 'lutff_global/s_r')
// (2, 9, 'neigh_op_bnl_0')
// (2, 11, 'lutff_global/s_r')
// (6, 8, 'lutff_global/s_r')
// (6, 14, 'lutff_global/s_r')

reg n5 = 0;
// (0, 0, 'glb_netwk_7')
// (2, 2, 'glb2local_1')
// (2, 2, 'local_g0_5')
// (2, 2, 'lutff_4/in_3')
// (4, 3, 'glb2local_0')
// (4, 3, 'glb2local_1')
// (4, 3, 'local_g0_4')
// (4, 3, 'local_g0_5')
// (4, 3, 'lutff_1/in_3')
// (4, 3, 'lutff_2/in_3')
// (5, 2, 'glb2local_0')
// (5, 2, 'glb2local_3')
// (5, 2, 'local_g0_4')
// (5, 2, 'local_g0_7')
// (5, 2, 'lutff_1/in_3')
// (5, 2, 'lutff_2/in_3')
// (5, 3, 'glb2local_0')
// (5, 3, 'local_g0_4')
// (5, 3, 'lutff_5/in_3')
// (6, 4, 'glb2local_1')
// (6, 4, 'local_g0_5')
// (6, 4, 'lutff_4/in_3')
// (8, 5, 'lutff_global/cen')
// (8, 5, 'neigh_op_tnr_1')
// (8, 5, 'sp4_r_v_b_47')
// (8, 6, 'lutff_global/cen')
// (8, 6, 'neigh_op_rgt_1')
// (8, 6, 'sp4_r_v_b_34')
// (8, 7, 'lutff_global/cen')
// (8, 7, 'neigh_op_bnr_1')
// (8, 7, 'sp4_r_v_b_23')
// (8, 8, 'lutff_global/cen')
// (8, 8, 'sp4_r_v_b_10')
// (9, 4, 'glb2local_2')
// (9, 4, 'local_g0_6')
// (9, 4, 'lutff_4/in_2')
// (9, 4, 'sp4_v_t_47')
// (9, 5, 'neigh_op_top_1')
// (9, 5, 'sp4_v_b_47')
// (9, 6, 'lutff_1/out')
// (9, 6, 'sp4_v_b_34')
// (9, 7, 'neigh_op_bot_1')
// (9, 7, 'sp4_v_b_23')
// (9, 8, 'sp4_h_r_4')
// (9, 8, 'sp4_v_b_10')
// (10, 5, 'neigh_op_tnl_1')
// (10, 6, 'neigh_op_lft_1')
// (10, 7, 'neigh_op_bnl_1')
// (10, 8, 'sp4_h_r_17')
// (11, 4, 'glb2local_0')
// (11, 4, 'local_g0_4')
// (11, 4, 'lutff_6/in_0')
// (11, 6, 'lutff_global/cen')
// (11, 8, 'sp4_h_r_28')
// (12, 8, 'sp4_h_r_41')
// (13, 8, 'fabout')
// (13, 8, 'local_g0_1')
// (13, 8, 'span4_horz_41')

wire n6;
// (0, 2, 'span12_horz_0')
// (1, 2, 'sp12_h_r_3')
// (2, 2, 'local_g0_4')
// (2, 2, 'lutff_4/in_2')
// (2, 2, 'sp12_h_r_4')
// (3, 1, 'neigh_op_tnr_0')
// (3, 2, 'neigh_op_rgt_0')
// (3, 2, 'sp12_h_r_7')
// (3, 3, 'neigh_op_bnr_0')
// (4, 1, 'neigh_op_top_0')
// (4, 2, 'lutff_0/out')
// (4, 2, 'sp12_h_r_8')
// (4, 3, 'neigh_op_bot_0')
// (5, 1, 'neigh_op_tnl_0')
// (5, 2, 'local_g1_0')
// (5, 2, 'lutff_7/in_0')
// (5, 2, 'neigh_op_lft_0')
// (5, 2, 'sp12_h_r_11')
// (5, 3, 'neigh_op_bnl_0')
// (6, 2, 'sp12_h_r_12')
// (7, 2, 'sp12_h_r_15')
// (8, 2, 'sp12_h_r_16')
// (9, 2, 'sp12_h_r_19')
// (10, 2, 'sp12_h_r_20')
// (11, 2, 'sp12_h_r_23')
// (12, 2, 'sp12_h_l_23')

wire n7;
// (0, 2, 'span12_horz_5')
// (1, 2, 'sp12_h_r_6')
// (2, 2, 'local_g0_1')
// (2, 2, 'lutff_0/in_1')
// (2, 2, 'sp12_h_r_9')
// (3, 2, 'sp12_h_r_10')
// (4, 1, 'neigh_op_tnr_3')
// (4, 2, 'neigh_op_rgt_3')
// (4, 2, 'sp12_h_r_13')
// (4, 3, 'neigh_op_bnr_3')
// (5, 1, 'neigh_op_top_3')
// (5, 2, 'local_g0_3')
// (5, 2, 'local_g1_3')
// (5, 2, 'lutff_2/in_2')
// (5, 2, 'lutff_3/out')
// (5, 2, 'lutff_6/in_1')
// (5, 2, 'sp12_h_r_14')
// (5, 3, 'neigh_op_bot_3')
// (6, 1, 'neigh_op_tnl_3')
// (6, 2, 'neigh_op_lft_3')
// (6, 2, 'sp12_h_r_17')
// (6, 3, 'neigh_op_bnl_3')
// (7, 2, 'sp12_h_r_18')
// (8, 2, 'sp12_h_r_21')
// (9, 2, 'sp12_h_r_22')
// (10, 2, 'sp12_h_l_22')

wire n8;
// (0, 3, 'span12_horz_10')
// (1, 3, 'sp12_h_r_13')
// (2, 3, 'sp12_h_r_14')
// (3, 3, 'sp12_h_r_17')
// (4, 3, 'local_g0_2')
// (4, 3, 'lutff_7/in_1')
// (4, 3, 'sp12_h_r_18')
// (5, 2, 'neigh_op_tnr_7')
// (5, 3, 'local_g3_7')
// (5, 3, 'lutff_6/in_0')
// (5, 3, 'neigh_op_rgt_7')
// (5, 3, 'sp12_h_r_21')
// (5, 4, 'neigh_op_bnr_7')
// (6, 2, 'neigh_op_top_7')
// (6, 3, 'lutff_7/out')
// (6, 3, 'sp12_h_r_22')
// (6, 4, 'neigh_op_bot_7')
// (7, 2, 'neigh_op_tnl_7')
// (7, 3, 'local_g0_7')
// (7, 3, 'local_g1_7')
// (7, 3, 'lutff_1/in_3')
// (7, 3, 'lutff_7/in_0')
// (7, 3, 'neigh_op_lft_7')
// (7, 3, 'sp12_h_l_22')
// (7, 4, 'neigh_op_bnl_7')

reg n9 = 0;
// (0, 3, 'span12_horz_12')
// (0, 3, 'span4_horz_0')
// (1, 2, 'neigh_op_tnr_4')
// (1, 3, 'neigh_op_rgt_4')
// (1, 3, 'sp12_h_r_15')
// (1, 3, 'sp4_h_r_13')
// (1, 3, 'sp4_h_r_9')
// (1, 4, 'neigh_op_bnr_4')
// (2, 2, 'local_g1_4')
// (2, 2, 'lutff_0/in_3')
// (2, 2, 'neigh_op_top_4')
// (2, 3, 'local_g0_4')
// (2, 3, 'lutff_4/in_2')
// (2, 3, 'lutff_4/out')
// (2, 3, 'sp12_h_r_16')
// (2, 3, 'sp4_h_r_20')
// (2, 3, 'sp4_h_r_24')
// (2, 3, 'sp4_h_r_8')
// (2, 4, 'neigh_op_bot_4')
// (3, 1, 'sp4_r_v_b_30')
// (3, 2, 'neigh_op_tnl_4')
// (3, 2, 'sp4_r_v_b_19')
// (3, 3, 'neigh_op_lft_4')
// (3, 3, 'sp12_h_r_19')
// (3, 3, 'sp4_h_r_21')
// (3, 3, 'sp4_h_r_33')
// (3, 3, 'sp4_h_r_37')
// (3, 3, 'sp4_r_v_b_6')
// (3, 4, 'neigh_op_bnl_4')
// (4, 0, 'span4_vert_30')
// (4, 1, 'sp4_r_v_b_27')
// (4, 1, 'sp4_v_b_30')
// (4, 2, 'local_g0_3')
// (4, 2, 'lutff_0/in_3')
// (4, 2, 'sp4_r_v_b_14')
// (4, 2, 'sp4_v_b_19')
// (4, 3, 'local_g1_4')
// (4, 3, 'local_g2_0')
// (4, 3, 'lutff_1/in_2')
// (4, 3, 'lutff_2/in_0')
// (4, 3, 'sp12_h_r_20')
// (4, 3, 'sp4_h_l_37')
// (4, 3, 'sp4_h_r_32')
// (4, 3, 'sp4_h_r_44')
// (4, 3, 'sp4_r_v_b_3')
// (4, 3, 'sp4_v_b_6')
// (5, 0, 'span4_vert_27')
// (5, 1, 'sp4_v_b_27')
// (5, 2, 'local_g0_6')
// (5, 2, 'local_g1_6')
// (5, 2, 'lutff_1/in_1')
// (5, 2, 'lutff_2/in_1')
// (5, 2, 'sp4_v_b_14')
// (5, 3, 'local_g0_7')
// (5, 3, 'local_g1_7')
// (5, 3, 'lutff_0/in_1')
// (5, 3, 'lutff_1/in_3')
// (5, 3, 'lutff_3/in_0')
// (5, 3, 'sp12_h_r_23')
// (5, 3, 'sp4_h_l_44')
// (5, 3, 'sp4_h_r_45')
// (5, 3, 'sp4_v_b_3')
// (6, 3, 'sp12_h_l_23')
// (6, 3, 'sp4_h_l_45')

reg n10 = 0;
// (0, 3, 'span12_horz_14')
// (1, 2, 'neigh_op_tnr_5')
// (1, 3, 'neigh_op_rgt_5')
// (1, 3, 'sp12_h_r_17')
// (1, 4, 'neigh_op_bnr_5')
// (2, 2, 'neigh_op_top_5')
// (2, 3, 'local_g0_5')
// (2, 3, 'lutff_5/in_2')
// (2, 3, 'lutff_5/out')
// (2, 3, 'sp12_h_r_18')
// (2, 4, 'neigh_op_bot_5')
// (3, 2, 'neigh_op_tnl_5')
// (3, 3, 'neigh_op_lft_5')
// (3, 3, 'sp12_h_r_21')
// (3, 3, 'sp4_h_r_10')
// (3, 4, 'neigh_op_bnl_5')
// (4, 1, 'sp4_r_v_b_36')
// (4, 2, 'local_g1_1')
// (4, 2, 'lutff_0/in_2')
// (4, 2, 'sp4_r_v_b_25')
// (4, 3, 'local_g0_6')
// (4, 3, 'local_g1_6')
// (4, 3, 'lutff_1/in_1')
// (4, 3, 'lutff_2/in_1')
// (4, 3, 'sp12_h_r_22')
// (4, 3, 'sp4_h_r_23')
// (4, 3, 'sp4_r_v_b_12')
// (4, 4, 'sp4_r_v_b_1')
// (5, 0, 'span12_vert_5')
// (5, 0, 'span4_vert_36')
// (5, 1, 'sp12_v_b_5')
// (5, 1, 'sp4_v_b_36')
// (5, 2, 'local_g2_2')
// (5, 2, 'local_g3_2')
// (5, 2, 'lutff_3/in_3')
// (5, 2, 'lutff_4/in_1')
// (5, 2, 'sp12_v_b_2')
// (5, 2, 'sp4_v_b_25')
// (5, 3, 'local_g1_4')
// (5, 3, 'local_g2_2')
// (5, 3, 'lutff_0/in_3')
// (5, 3, 'lutff_1/in_1')
// (5, 3, 'lutff_5/in_2')
// (5, 3, 'sp12_h_l_22')
// (5, 3, 'sp12_v_b_1')
// (5, 3, 'sp4_h_r_34')
// (5, 3, 'sp4_v_b_12')
// (5, 4, 'sp4_v_b_1')
// (6, 3, 'sp4_h_r_47')
// (7, 3, 'sp4_h_l_47')

reg n11 = 0;
// (0, 3, 'span12_horz_2')
// (1, 2, 'neigh_op_tnr_7')
// (1, 3, 'neigh_op_rgt_7')
// (1, 3, 'sp12_h_r_5')
// (1, 3, 'sp4_h_r_2')
// (1, 4, 'neigh_op_bnr_7')
// (2, 2, 'local_g0_7')
// (2, 2, 'local_g1_7')
// (2, 2, 'lutff_0/in_2')
// (2, 2, 'lutff_4/in_1')
// (2, 2, 'neigh_op_top_7')
// (2, 3, 'local_g2_7')
// (2, 3, 'lutff_7/in_2')
// (2, 3, 'lutff_7/out')
// (2, 3, 'sp12_h_r_6')
// (2, 3, 'sp4_h_r_15')
// (2, 4, 'neigh_op_bot_7')
// (3, 2, 'neigh_op_tnl_7')
// (3, 3, 'neigh_op_lft_7')
// (3, 3, 'sp12_h_r_9')
// (3, 3, 'sp4_h_r_26')
// (3, 4, 'neigh_op_bnl_7')
// (4, 1, 'sp4_r_v_b_32')
// (4, 2, 'sp4_r_v_b_21')
// (4, 3, 'local_g1_2')
// (4, 3, 'lutff_5/in_2')
// (4, 3, 'sp12_h_r_10')
// (4, 3, 'sp4_h_r_39')
// (4, 3, 'sp4_r_v_b_8')
// (5, 0, 'span4_vert_32')
// (5, 1, 'sp4_v_b_32')
// (5, 2, 'local_g0_5')
// (5, 2, 'local_g1_5')
// (5, 2, 'lutff_1/in_2')
// (5, 2, 'lutff_2/in_0')
// (5, 2, 'lutff_4/in_0')
// (5, 2, 'sp4_v_b_21')
// (5, 3, 'local_g0_6')
// (5, 3, 'local_g1_6')
// (5, 3, 'lutff_0/in_2')
// (5, 3, 'lutff_1/in_2')
// (5, 3, 'lutff_3/in_1')
// (5, 3, 'sp12_h_r_13')
// (5, 3, 'sp4_h_l_39')
// (5, 3, 'sp4_h_r_6')
// (5, 3, 'sp4_v_b_8')
// (6, 3, 'sp12_h_r_14')
// (6, 3, 'sp4_h_r_19')
// (7, 3, 'sp12_h_r_17')
// (7, 3, 'sp4_h_r_30')
// (8, 3, 'sp12_h_r_18')
// (8, 3, 'sp4_h_r_43')
// (9, 3, 'sp12_h_r_21')
// (9, 3, 'sp4_h_l_43')
// (10, 3, 'sp12_h_r_22')
// (11, 3, 'sp12_h_l_22')

wire n12;
// (0, 3, 'span12_horz_7')
// (1, 3, 'sp12_h_r_8')
// (2, 3, 'sp12_h_r_11')
// (3, 3, 'sp12_h_r_12')
// (4, 3, 'sp12_h_r_15')
// (5, 3, 'sp12_h_r_16')
// (6, 2, 'local_g3_6')
// (6, 2, 'lutff_2/in_1')
// (6, 2, 'neigh_op_tnr_6')
// (6, 3, 'local_g0_3')
// (6, 3, 'lutff_4/in_3')
// (6, 3, 'neigh_op_rgt_6')
// (6, 3, 'sp12_h_r_19')
// (6, 4, 'neigh_op_bnr_6')
// (7, 2, 'neigh_op_top_6')
// (7, 3, 'lutff_6/out')
// (7, 3, 'sp12_h_r_20')
// (7, 4, 'neigh_op_bot_6')
// (8, 2, 'neigh_op_tnl_6')
// (8, 3, 'neigh_op_lft_6')
// (8, 3, 'sp12_h_r_23')
// (8, 4, 'neigh_op_bnl_6')
// (9, 3, 'sp12_h_l_23')

reg n13 = 0;
// (0, 4, 'span12_horz_1')
// (1, 4, 'sp12_h_r_2')
// (2, 4, 'sp12_h_r_5')
// (3, 4, 'sp12_h_r_6')
// (4, 4, 'sp12_h_r_9')
// (5, 4, 'sp12_h_r_10')
// (5, 6, 'sp4_h_r_7')
// (6, 4, 'sp12_h_r_13')
// (6, 6, 'sp4_h_r_18')
// (7, 4, 'sp12_h_r_14')
// (7, 6, 'sp4_h_r_31')
// (8, 3, 'neigh_op_tnr_5')
// (8, 3, 'sp4_r_v_b_39')
// (8, 4, 'neigh_op_rgt_5')
// (8, 4, 'sp12_h_r_17')
// (8, 4, 'sp4_r_v_b_26')
// (8, 5, 'local_g0_5')
// (8, 5, 'local_g1_5')
// (8, 5, 'lutff_0/in_2')
// (8, 5, 'lutff_1/in_2')
// (8, 5, 'lutff_3/in_2')
// (8, 5, 'neigh_op_bnr_5')
// (8, 5, 'sp4_r_v_b_15')
// (8, 6, 'local_g1_2')
// (8, 6, 'local_g2_2')
// (8, 6, 'lutff_0/in_2')
// (8, 6, 'lutff_1/in_2')
// (8, 6, 'lutff_2/in_2')
// (8, 6, 'lutff_3/in_2')
// (8, 6, 'lutff_4/in_2')
// (8, 6, 'sp4_h_r_42')
// (8, 6, 'sp4_r_v_b_2')
// (8, 7, 'local_g2_5')
// (8, 7, 'local_g3_7')
// (8, 7, 'lutff_0/in_3')
// (8, 7, 'lutff_1/in_2')
// (8, 7, 'lutff_3/in_2')
// (8, 7, 'lutff_4/in_2')
// (8, 7, 'sp4_r_v_b_37')
// (8, 7, 'sp4_r_v_b_47')
// (8, 8, 'sp4_r_v_b_24')
// (8, 8, 'sp4_r_v_b_34')
// (8, 9, 'sp4_r_v_b_13')
// (8, 9, 'sp4_r_v_b_23')
// (8, 10, 'sp4_r_v_b_0')
// (8, 10, 'sp4_r_v_b_10')
// (9, 2, 'sp4_v_t_39')
// (9, 3, 'neigh_op_top_5')
// (9, 3, 'sp4_v_b_39')
// (9, 4, 'local_g2_5')
// (9, 4, 'local_g3_5')
// (9, 4, 'lutff_0/in_3')
// (9, 4, 'lutff_1/in_2')
// (9, 4, 'lutff_5/in_1')
// (9, 4, 'lutff_5/out')
// (9, 4, 'sp12_h_r_18')
// (9, 4, 'sp4_v_b_26')
// (9, 5, 'neigh_op_bot_5')
// (9, 5, 'sp4_v_b_15')
// (9, 6, 'sp4_h_l_42')
// (9, 6, 'sp4_h_r_0')
// (9, 6, 'sp4_v_b_2')
// (9, 6, 'sp4_v_t_37')
// (9, 6, 'sp4_v_t_47')
// (9, 7, 'sp4_v_b_37')
// (9, 7, 'sp4_v_b_47')
// (9, 8, 'sp4_v_b_24')
// (9, 8, 'sp4_v_b_34')
// (9, 9, 'sp4_v_b_13')
// (9, 9, 'sp4_v_b_23')
// (9, 10, 'sp4_v_b_0')
// (9, 10, 'sp4_v_b_10')
// (10, 3, 'neigh_op_tnl_5')
// (10, 4, 'neigh_op_lft_5')
// (10, 4, 'sp12_h_r_21')
// (10, 5, 'neigh_op_bnl_5')
// (10, 6, 'sp4_h_r_13')
// (11, 4, 'local_g0_6')
// (11, 4, 'lutff_5/in_3')
// (11, 4, 'lutff_6/in_2')
// (11, 4, 'lutff_7/in_1')
// (11, 4, 'sp12_h_r_22')
// (11, 6, 'local_g2_0')
// (11, 6, 'lutff_2/in_2')
// (11, 6, 'lutff_4/in_2')
// (11, 6, 'sp4_h_r_24')
// (12, 4, 'sp12_h_l_22')
// (12, 6, 'sp4_h_r_37')
// (13, 6, 'span4_horz_37')

wire n14;
// (0, 4, 'span4_horz_1')
// (0, 10, 'span12_horz_3')
// (1, 4, 'sp12_h_r_0')
// (1, 4, 'sp4_h_r_12')
// (1, 10, 'sp12_h_r_4')
// (2, 4, 'sp12_h_r_3')
// (2, 4, 'sp4_h_r_25')
// (2, 10, 'sp12_h_r_7')
// (3, 4, 'sp12_h_r_4')
// (3, 4, 'sp4_h_r_36')
// (3, 5, 'sp4_r_v_b_36')
// (3, 6, 'sp4_r_v_b_25')
// (3, 7, 'sp4_r_v_b_12')
// (3, 8, 'sp4_r_v_b_1')
// (3, 10, 'sp12_h_r_8')
// (4, 4, 'sp12_h_r_7')
// (4, 4, 'sp4_h_l_36')
// (4, 4, 'sp4_v_t_36')
// (4, 5, 'local_g2_4')
// (4, 5, 'lutff_4/in_0')
// (4, 5, 'lutff_7/in_1')
// (4, 5, 'sp4_v_b_36')
// (4, 6, 'sp4_v_b_25')
// (4, 7, 'sp4_v_b_12')
// (4, 8, 'sp4_h_r_7')
// (4, 8, 'sp4_v_b_1')
// (4, 10, 'sp12_h_r_11')
// (5, 4, 'local_g1_0')
// (5, 4, 'lutff_6/in_1')
// (5, 4, 'sp12_h_r_8')
// (5, 8, 'sp4_h_r_18')
// (5, 10, 'local_g0_4')
// (5, 10, 'lutff_1/in_1')
// (5, 10, 'sp12_h_r_12')
// (6, 4, 'sp12_h_r_11')
// (6, 8, 'sp4_h_r_31')
// (6, 10, 'sp12_h_r_15')
// (7, 4, 'sp12_h_r_12')
// (7, 8, 'sp4_h_r_42')
// (7, 9, 'sp4_r_v_b_37')
// (7, 10, 'sp12_h_r_16')
// (7, 10, 'sp4_r_v_b_24')
// (7, 11, 'sp4_r_v_b_13')
// (7, 12, 'sp4_r_v_b_0')
// (8, 4, 'sp12_h_r_15')
// (8, 8, 'sp4_h_l_42')
// (8, 8, 'sp4_v_t_37')
// (8, 9, 'sp4_v_b_37')
// (8, 10, 'sp12_h_r_19')
// (8, 10, 'sp4_v_b_24')
// (8, 11, 'local_g0_5')
// (8, 11, 'lutff_2/in_1')
// (8, 11, 'sp4_v_b_13')
// (8, 12, 'sp4_v_b_0')
// (9, 4, 'sp12_h_r_0')
// (9, 4, 'sp12_h_r_16')
// (9, 4, 'sp12_v_t_23')
// (9, 5, 'sp12_v_b_23')
// (9, 6, 'sp12_v_b_20')
// (9, 7, 'sp12_v_b_19')
// (9, 8, 'sp12_v_b_16')
// (9, 9, 'local_g2_7')
// (9, 9, 'local_g3_7')
// (9, 9, 'lutff_1/in_1')
// (9, 9, 'lutff_7/in_0')
// (9, 9, 'sp12_v_b_15')
// (9, 10, 'sp12_h_r_20')
// (9, 10, 'sp12_v_b_12')
// (9, 11, 'sp12_v_b_11')
// (9, 12, 'sp12_v_b_8')
// (9, 13, 'sp12_v_b_7')
// (9, 14, 'sp12_v_b_4')
// (9, 15, 'sp12_v_b_3')
// (9, 16, 'sp12_v_b_0')
// (10, 3, 'neigh_op_tnr_6')
// (10, 4, 'neigh_op_rgt_6')
// (10, 4, 'sp12_h_r_19')
// (10, 4, 'sp12_h_r_3')
// (10, 5, 'neigh_op_bnr_6')
// (10, 10, 'sp12_h_r_23')
// (11, 0, 'span12_vert_19')
// (11, 1, 'sp12_v_b_19')
// (11, 2, 'sp12_v_b_16')
// (11, 3, 'neigh_op_top_6')
// (11, 3, 'sp12_v_b_15')
// (11, 4, 'lutff_6/out')
// (11, 4, 'sp12_h_r_20')
// (11, 4, 'sp12_h_r_4')
// (11, 4, 'sp12_v_b_12')
// (11, 5, 'neigh_op_bot_6')
// (11, 5, 'sp12_v_b_11')
// (11, 6, 'sp12_v_b_8')
// (11, 7, 'sp12_v_b_7')
// (11, 8, 'local_g2_4')
// (11, 8, 'lutff_1/in_3')
// (11, 8, 'sp12_v_b_4')
// (11, 9, 'sp12_v_b_3')
// (11, 10, 'sp12_h_l_23')
// (11, 10, 'sp12_v_b_0')
// (11, 10, 'sp12_v_t_23')
// (11, 11, 'local_g3_7')
// (11, 11, 'lutff_5/in_1')
// (11, 11, 'sp12_v_b_23')
// (11, 12, 'sp12_v_b_20')
// (11, 13, 'sp12_v_b_19')
// (11, 14, 'sp12_v_b_16')
// (11, 15, 'sp12_v_b_15')
// (11, 16, 'sp12_v_b_12')
// (11, 17, 'span12_vert_11')
// (12, 3, 'neigh_op_tnl_6')
// (12, 4, 'neigh_op_lft_6')
// (12, 4, 'sp12_h_r_23')
// (12, 4, 'sp12_h_r_7')
// (12, 5, 'neigh_op_bnl_6')
// (13, 4, 'span12_horz_23')
// (13, 4, 'span12_horz_7')

reg n15 = 0;
// (0, 5, 'span12_horz_10')
// (1, 4, 'neigh_op_tnr_3')
// (1, 5, 'neigh_op_rgt_3')
// (1, 5, 'sp12_h_r_13')
// (1, 6, 'neigh_op_bnr_3')
// (1, 12, 'sp4_r_v_b_38')
// (1, 13, 'sp4_r_v_b_27')
// (1, 14, 'sp4_r_v_b_14')
// (1, 14, 'sp4_r_v_b_36')
// (1, 15, 'sp4_r_v_b_25')
// (1, 15, 'sp4_r_v_b_3')
// (1, 16, 'sp4_r_v_b_12')
// (2, 4, 'neigh_op_top_3')
// (2, 4, 'sp12_v_t_22')
// (2, 5, 'lutff_3/out')
// (2, 5, 'sp12_h_r_14')
// (2, 5, 'sp12_v_b_22')
// (2, 6, 'neigh_op_bot_3')
// (2, 6, 'sp12_v_b_21')
// (2, 7, 'sp12_v_b_18')
// (2, 8, 'sp12_v_b_17')
// (2, 9, 'sp12_v_b_14')
// (2, 10, 'sp12_v_b_13')
// (2, 11, 'sp12_v_b_10')
// (2, 11, 'sp4_h_r_8')
// (2, 11, 'sp4_v_t_38')
// (2, 12, 'local_g2_1')
// (2, 12, 'lutff_0/in_3')
// (2, 12, 'sp12_v_b_9')
// (2, 12, 'sp4_v_b_38')
// (2, 13, 'sp12_v_b_6')
// (2, 13, 'sp4_h_r_1')
// (2, 13, 'sp4_v_b_27')
// (2, 13, 'sp4_v_t_36')
// (2, 14, 'sp12_v_b_5')
// (2, 14, 'sp4_v_b_14')
// (2, 14, 'sp4_v_b_36')
// (2, 15, 'sp12_v_b_2')
// (2, 15, 'sp4_v_b_25')
// (2, 15, 'sp4_v_b_3')
// (2, 16, 'sp12_v_b_1')
// (2, 16, 'sp4_v_b_12')
// (2, 17, 'span4_vert_1')
// (3, 4, 'neigh_op_tnl_3')
// (3, 5, 'neigh_op_lft_3')
// (3, 5, 'sp12_h_r_17')
// (3, 6, 'neigh_op_bnl_3')
// (3, 10, 'sp4_h_r_5')
// (3, 11, 'sp4_h_r_21')
// (3, 12, 'sp4_h_r_7')
// (3, 13, 'sp4_h_r_12')
// (3, 14, 'sp4_h_r_5')
// (4, 5, 'sp12_h_r_18')
// (4, 10, 'local_g0_0')
// (4, 10, 'lutff_0/in_2')
// (4, 10, 'sp4_h_r_16')
// (4, 11, 'local_g2_0')
// (4, 11, 'lutff_0/in_2')
// (4, 11, 'lutff_1/in_1')
// (4, 11, 'sp4_h_r_32')
// (4, 12, 'local_g0_2')
// (4, 12, 'lutff_6/in_2')
// (4, 12, 'sp4_h_r_18')
// (4, 13, 'local_g2_1')
// (4, 13, 'lutff_5/in_2')
// (4, 13, 'sp4_h_r_25')
// (4, 14, 'local_g0_0')
// (4, 14, 'lutff_6/in_2')
// (4, 14, 'sp4_h_r_16')
// (5, 4, 'sp4_r_v_b_41')
// (5, 5, 'sp12_h_r_21')
// (5, 5, 'sp4_h_r_10')
// (5, 5, 'sp4_r_v_b_28')
// (5, 6, 'sp4_r_v_b_17')
// (5, 7, 'local_g1_4')
// (5, 7, 'lutff_4/in_3')
// (5, 7, 'sp4_r_v_b_4')
// (5, 8, 'sp4_r_v_b_36')
// (5, 9, 'sp4_r_v_b_25')
// (5, 10, 'sp4_h_r_29')
// (5, 10, 'sp4_r_v_b_12')
// (5, 11, 'sp4_h_r_45')
// (5, 11, 'sp4_r_v_b_1')
// (5, 12, 'local_g2_4')
// (5, 12, 'lutff_0/in_2')
// (5, 12, 'lutff_1/in_1')
// (5, 12, 'lutff_3/in_1')
// (5, 12, 'sp4_h_r_31')
// (5, 12, 'sp4_r_v_b_36')
// (5, 12, 'sp4_r_v_b_45')
// (5, 13, 'local_g0_3')
// (5, 13, 'local_g1_1')
// (5, 13, 'lutff_0/in_2')
// (5, 13, 'lutff_2/in_3')
// (5, 13, 'sp4_h_r_36')
// (5, 13, 'sp4_r_v_b_25')
// (5, 13, 'sp4_r_v_b_32')
// (5, 14, 'local_g2_4')
// (5, 14, 'lutff_5/in_3')
// (5, 14, 'sp4_h_r_29')
// (5, 14, 'sp4_r_v_b_12')
// (5, 14, 'sp4_r_v_b_21')
// (5, 15, 'sp4_r_v_b_1')
// (5, 15, 'sp4_r_v_b_8')
// (6, 3, 'sp4_v_t_41')
// (6, 4, 'sp4_v_b_41')
// (6, 5, 'sp12_h_r_22')
// (6, 5, 'sp4_h_r_23')
// (6, 5, 'sp4_v_b_28')
// (6, 6, 'sp4_v_b_17')
// (6, 7, 'local_g1_4')
// (6, 7, 'lutff_1/in_2')
// (6, 7, 'lutff_4/in_1')
// (6, 7, 'sp4_h_r_1')
// (6, 7, 'sp4_v_b_4')
// (6, 7, 'sp4_v_t_36')
// (6, 8, 'local_g2_4')
// (6, 8, 'lutff_1/in_1')
// (6, 8, 'sp4_v_b_36')
// (6, 9, 'local_g3_1')
// (6, 9, 'lutff_0/in_2')
// (6, 9, 'sp4_r_v_b_42')
// (6, 9, 'sp4_v_b_25')
// (6, 10, 'local_g1_4')
// (6, 10, 'lutff_4/in_3')
// (6, 10, 'sp4_h_r_40')
// (6, 10, 'sp4_r_v_b_31')
// (6, 10, 'sp4_v_b_12')
// (6, 11, 'sp4_h_l_45')
// (6, 11, 'sp4_r_v_b_18')
// (6, 11, 'sp4_r_v_b_40')
// (6, 11, 'sp4_v_b_1')
// (6, 11, 'sp4_v_t_36')
// (6, 11, 'sp4_v_t_45')
// (6, 12, 'local_g2_4')
// (6, 12, 'lutff_4/in_2')
// (6, 12, 'sp4_h_r_42')
// (6, 12, 'sp4_r_v_b_29')
// (6, 12, 'sp4_r_v_b_7')
// (6, 12, 'sp4_v_b_36')
// (6, 12, 'sp4_v_b_45')
// (6, 13, 'sp4_h_l_36')
// (6, 13, 'sp4_h_r_1')
// (6, 13, 'sp4_r_v_b_16')
// (6, 13, 'sp4_v_b_25')
// (6, 13, 'sp4_v_b_32')
// (6, 14, 'sp4_h_r_40')
// (6, 14, 'sp4_r_v_b_5')
// (6, 14, 'sp4_v_b_12')
// (6, 14, 'sp4_v_b_21')
// (6, 15, 'sp4_v_b_1')
// (6, 15, 'sp4_v_b_8')
// (7, 5, 'sp12_h_l_22')
// (7, 5, 'sp12_v_t_22')
// (7, 5, 'sp4_h_r_34')
// (7, 6, 'sp12_v_b_22')
// (7, 7, 'local_g0_4')
// (7, 7, 'lutff_6/in_2')
// (7, 7, 'sp12_v_b_21')
// (7, 7, 'sp4_h_r_12')
// (7, 8, 'sp12_v_b_18')
// (7, 8, 'sp4_v_t_42')
// (7, 9, 'sp12_v_b_17')
// (7, 9, 'sp4_v_b_42')
// (7, 10, 'sp12_v_b_14')
// (7, 10, 'sp4_h_l_40')
// (7, 10, 'sp4_h_r_8')
// (7, 10, 'sp4_v_b_31')
// (7, 10, 'sp4_v_t_40')
// (7, 11, 'sp12_v_b_13')
// (7, 11, 'sp4_v_b_18')
// (7, 11, 'sp4_v_b_40')
// (7, 12, 'sp12_v_b_10')
// (7, 12, 'sp4_h_l_42')
// (7, 12, 'sp4_h_r_10')
// (7, 12, 'sp4_v_b_29')
// (7, 12, 'sp4_v_b_7')
// (7, 13, 'local_g0_4')
// (7, 13, 'local_g1_4')
// (7, 13, 'lutff_0/in_2')
// (7, 13, 'lutff_1/in_1')
// (7, 13, 'lutff_6/in_3')
// (7, 13, 'sp12_v_b_9')
// (7, 13, 'sp4_h_r_12')
// (7, 13, 'sp4_v_b_16')
// (7, 14, 'local_g3_6')
// (7, 14, 'lutff_5/in_2')
// (7, 14, 'sp12_v_b_6')
// (7, 14, 'sp4_h_l_40')
// (7, 14, 'sp4_v_b_5')
// (7, 15, 'sp12_v_b_5')
// (7, 16, 'sp12_v_b_2')
// (7, 17, 'span12_vert_1')
// (8, 5, 'sp4_h_r_47')
// (8, 6, 'sp4_r_v_b_38')
// (8, 7, 'sp4_h_r_25')
// (8, 7, 'sp4_r_v_b_27')
// (8, 8, 'sp4_r_v_b_14')
// (8, 9, 'local_g1_3')
// (8, 9, 'lutff_1/in_1')
// (8, 9, 'lutff_2/in_2')
// (8, 9, 'lutff_7/in_3')
// (8, 9, 'sp4_r_v_b_3')
// (8, 10, 'local_g0_5')
// (8, 10, 'lutff_1/in_2')
// (8, 10, 'sp4_h_r_21')
// (8, 12, 'local_g0_7')
// (8, 12, 'lutff_0/in_1')
// (8, 12, 'sp4_h_r_23')
// (8, 13, 'local_g2_1')
// (8, 13, 'lutff_1/in_2')
// (8, 13, 'lutff_5/in_2')
// (8, 13, 'lutff_6/in_3')
// (8, 13, 'sp4_h_r_25')
// (9, 5, 'sp4_h_l_47')
// (9, 5, 'sp4_v_t_38')
// (9, 6, 'sp4_v_b_38')
// (9, 7, 'sp4_h_r_36')
// (9, 7, 'sp4_v_b_27')
// (9, 8, 'sp4_v_b_14')
// (9, 9, 'sp4_v_b_3')
// (9, 10, 'sp4_h_r_32')
// (9, 12, 'sp4_h_r_34')
// (9, 13, 'sp4_h_r_36')
// (10, 7, 'sp4_h_l_36')
// (10, 10, 'sp4_h_r_45')
// (10, 12, 'sp4_h_r_47')
// (10, 13, 'sp4_h_l_36')
// (11, 10, 'sp4_h_l_45')
// (11, 12, 'sp4_h_l_47')

wire n16;
// (0, 5, 'span12_horz_13')
// (1, 5, 'sp12_h_r_14')
// (2, 5, 'sp12_h_r_17')
// (3, 5, 'sp12_h_r_18')
// (4, 5, 'sp12_h_r_21')
// (5, 5, 'local_g1_6')
// (5, 5, 'lutff_2/in_1')
// (5, 5, 'lutff_4/in_3')
// (5, 5, 'neigh_op_tnr_3')
// (5, 5, 'sp12_h_r_22')
// (5, 6, 'neigh_op_rgt_3')
// (5, 7, 'neigh_op_bnr_3')
// (6, 5, 'neigh_op_top_3')
// (6, 5, 'sp12_h_l_22')
// (6, 5, 'sp12_v_t_22')
// (6, 6, 'lutff_3/out')
// (6, 6, 'sp12_v_b_22')
// (6, 7, 'neigh_op_bot_3')
// (6, 7, 'sp12_v_b_21')
// (6, 8, 'sp12_v_b_18')
// (6, 9, 'sp12_v_b_17')
// (6, 10, 'sp12_v_b_14')
// (6, 11, 'sp12_v_b_13')
// (6, 12, 'sp12_v_b_10')
// (6, 13, 'sp12_v_b_9')
// (6, 14, 'sp12_v_b_6')
// (6, 15, 'sp12_v_b_5')
// (6, 16, 'sp12_v_b_2')
// (6, 17, 'span12_vert_1')
// (7, 5, 'local_g2_3')
// (7, 5, 'lutff_1/in_2')
// (7, 5, 'lutff_4/in_1')
// (7, 5, 'neigh_op_tnl_3')
// (7, 6, 'neigh_op_lft_3')
// (7, 7, 'neigh_op_bnl_3')

reg n17 = 0;
// (0, 5, 'span12_horz_4')
// (1, 5, 'sp12_h_r_7')
// (2, 5, 'sp12_h_r_8')
// (3, 4, 'neigh_op_tnr_2')
// (3, 5, 'neigh_op_rgt_2')
// (3, 5, 'sp12_h_r_11')
// (3, 6, 'neigh_op_bnr_2')
// (4, 4, 'neigh_op_top_2')
// (4, 5, 'local_g0_2')
// (4, 5, 'lutff_2/out')
// (4, 5, 'lutff_3/in_3')
// (4, 5, 'lutff_4/in_2')
// (4, 5, 'sp12_h_r_12')
// (4, 6, 'neigh_op_bot_2')
// (5, 4, 'neigh_op_tnl_2')
// (5, 5, 'local_g1_7')
// (5, 5, 'lutff_7/in_3')
// (5, 5, 'neigh_op_lft_2')
// (5, 5, 'sp12_h_r_15')
// (5, 6, 'neigh_op_bnl_2')
// (6, 5, 'sp12_h_r_16')
// (7, 5, 'sp12_h_r_19')
// (8, 5, 'sp12_h_r_20')
// (9, 5, 'sp12_h_r_23')
// (10, 5, 'sp12_h_l_23')

reg n18 = 0;
// (0, 5, 'span12_horz_8')
// (1, 4, 'neigh_op_tnr_2')
// (1, 5, 'neigh_op_rgt_2')
// (1, 5, 'sp12_h_r_11')
// (1, 6, 'neigh_op_bnr_2')
// (1, 10, 'sp4_r_v_b_39')
// (1, 11, 'sp4_r_v_b_26')
// (1, 12, 'sp4_r_v_b_15')
// (1, 12, 'sp4_r_v_b_37')
// (1, 13, 'sp4_r_v_b_2')
// (1, 13, 'sp4_r_v_b_24')
// (1, 14, 'sp4_r_v_b_13')
// (1, 15, 'sp4_r_v_b_0')
// (2, 3, 'sp12_v_t_23')
// (2, 4, 'neigh_op_top_2')
// (2, 4, 'sp12_v_b_23')
// (2, 5, 'lutff_2/out')
// (2, 5, 'sp12_h_r_12')
// (2, 5, 'sp12_v_b_20')
// (2, 6, 'neigh_op_bot_2')
// (2, 6, 'sp12_v_b_19')
// (2, 7, 'sp12_v_b_16')
// (2, 8, 'sp12_v_b_15')
// (2, 9, 'sp12_v_b_12')
// (2, 9, 'sp4_v_t_39')
// (2, 10, 'sp12_v_b_11')
// (2, 10, 'sp4_v_b_39')
// (2, 11, 'sp12_v_b_8')
// (2, 11, 'sp4_h_r_5')
// (2, 11, 'sp4_v_b_26')
// (2, 11, 'sp4_v_t_37')
// (2, 12, 'local_g3_7')
// (2, 12, 'lutff_0/in_2')
// (2, 12, 'sp12_v_b_7')
// (2, 12, 'sp4_v_b_15')
// (2, 12, 'sp4_v_b_37')
// (2, 13, 'sp12_v_b_4')
// (2, 13, 'sp4_h_r_8')
// (2, 13, 'sp4_v_b_2')
// (2, 13, 'sp4_v_b_24')
// (2, 14, 'sp12_v_b_3')
// (2, 14, 'sp4_v_b_13')
// (2, 15, 'sp12_v_b_0')
// (2, 15, 'sp4_v_b_0')
// (3, 4, 'neigh_op_tnl_2')
// (3, 5, 'neigh_op_lft_2')
// (3, 5, 'sp12_h_r_15')
// (3, 6, 'neigh_op_bnl_2')
// (3, 10, 'sp4_r_v_b_41')
// (3, 10, 'sp4_r_v_b_47')
// (3, 11, 'sp4_h_r_16')
// (3, 11, 'sp4_r_v_b_28')
// (3, 11, 'sp4_r_v_b_34')
// (3, 12, 'sp4_r_v_b_17')
// (3, 12, 'sp4_r_v_b_23')
// (3, 13, 'sp4_h_r_21')
// (3, 13, 'sp4_r_v_b_10')
// (3, 13, 'sp4_r_v_b_4')
// (3, 14, 'sp4_r_v_b_41')
// (3, 15, 'sp4_r_v_b_28')
// (3, 16, 'sp4_r_v_b_17')
// (4, 5, 'sp12_h_r_16')
// (4, 9, 'sp4_h_r_10')
// (4, 9, 'sp4_v_t_41')
// (4, 9, 'sp4_v_t_47')
// (4, 10, 'local_g2_1')
// (4, 10, 'lutff_0/in_3')
// (4, 10, 'sp4_v_b_41')
// (4, 10, 'sp4_v_b_47')
// (4, 11, 'local_g2_5')
// (4, 11, 'lutff_0/in_3')
// (4, 11, 'lutff_1/in_2')
// (4, 11, 'sp4_h_r_29')
// (4, 11, 'sp4_v_b_28')
// (4, 11, 'sp4_v_b_34')
// (4, 12, 'local_g0_7')
// (4, 12, 'lutff_6/in_3')
// (4, 12, 'sp4_v_b_17')
// (4, 12, 'sp4_v_b_23')
// (4, 13, 'local_g2_0')
// (4, 13, 'lutff_5/in_3')
// (4, 13, 'sp4_h_r_32')
// (4, 13, 'sp4_v_b_10')
// (4, 13, 'sp4_v_b_4')
// (4, 13, 'sp4_v_t_41')
// (4, 14, 'local_g2_1')
// (4, 14, 'lutff_6/in_3')
// (4, 14, 'sp4_v_b_41')
// (4, 15, 'sp4_v_b_28')
// (4, 16, 'sp4_v_b_17')
// (4, 17, 'span4_vert_4')
// (5, 4, 'sp4_r_v_b_45')
// (5, 5, 'sp12_h_r_19')
// (5, 5, 'sp4_r_v_b_32')
// (5, 6, 'sp4_r_v_b_21')
// (5, 7, 'local_g2_0')
// (5, 7, 'lutff_4/in_2')
// (5, 7, 'sp4_r_v_b_8')
// (5, 8, 'sp4_r_v_b_45')
// (5, 9, 'sp4_h_r_23')
// (5, 9, 'sp4_r_v_b_32')
// (5, 10, 'sp4_r_v_b_21')
// (5, 10, 'sp4_r_v_b_36')
// (5, 11, 'sp4_h_r_40')
// (5, 11, 'sp4_r_v_b_25')
// (5, 11, 'sp4_r_v_b_8')
// (5, 12, 'local_g3_0')
// (5, 12, 'lutff_0/in_3')
// (5, 12, 'lutff_1/in_2')
// (5, 12, 'lutff_3/in_2')
// (5, 12, 'sp4_r_v_b_12')
// (5, 12, 'sp4_r_v_b_40')
// (5, 13, 'local_g0_5')
// (5, 13, 'local_g1_5')
// (5, 13, 'lutff_0/in_3')
// (5, 13, 'lutff_2/in_2')
// (5, 13, 'sp4_h_r_45')
// (5, 13, 'sp4_r_v_b_1')
// (5, 13, 'sp4_r_v_b_29')
// (5, 14, 'local_g3_0')
// (5, 14, 'lutff_5/in_2')
// (5, 14, 'sp4_r_v_b_16')
// (5, 15, 'sp4_r_v_b_5')
// (6, 3, 'sp4_v_t_45')
// (6, 4, 'sp4_v_b_45')
// (6, 5, 'sp12_h_r_20')
// (6, 5, 'sp4_v_b_32')
// (6, 6, 'sp4_v_b_21')
// (6, 7, 'local_g0_0')
// (6, 7, 'local_g0_2')
// (6, 7, 'lutff_1/in_3')
// (6, 7, 'lutff_4/in_2')
// (6, 7, 'sp4_h_r_2')
// (6, 7, 'sp4_v_b_8')
// (6, 7, 'sp4_v_t_45')
// (6, 8, 'local_g2_5')
// (6, 8, 'lutff_1/in_2')
// (6, 8, 'sp4_v_b_45')
// (6, 9, 'local_g3_0')
// (6, 9, 'lutff_0/in_3')
// (6, 9, 'sp4_h_r_1')
// (6, 9, 'sp4_h_r_34')
// (6, 9, 'sp4_v_b_32')
// (6, 9, 'sp4_v_t_36')
// (6, 10, 'local_g1_5')
// (6, 10, 'lutff_4/in_2')
// (6, 10, 'sp4_v_b_21')
// (6, 10, 'sp4_v_b_36')
// (6, 11, 'sp4_h_l_40')
// (6, 11, 'sp4_v_b_25')
// (6, 11, 'sp4_v_b_8')
// (6, 11, 'sp4_v_t_40')
// (6, 12, 'local_g3_0')
// (6, 12, 'lutff_4/in_3')
// (6, 12, 'sp4_v_b_12')
// (6, 12, 'sp4_v_b_40')
// (6, 13, 'sp4_h_l_45')
// (6, 13, 'sp4_h_r_8')
// (6, 13, 'sp4_v_b_1')
// (6, 13, 'sp4_v_b_29')
// (6, 14, 'sp4_v_b_16')
// (6, 15, 'sp4_v_b_5')
// (7, 5, 'sp12_h_r_23')
// (7, 7, 'local_g0_7')
// (7, 7, 'lutff_6/in_3')
// (7, 7, 'sp4_h_r_15')
// (7, 9, 'sp4_h_r_12')
// (7, 9, 'sp4_h_r_47')
// (7, 10, 'sp4_r_v_b_41')
// (7, 11, 'sp4_r_v_b_28')
// (7, 12, 'sp4_r_v_b_17')
// (7, 13, 'local_g0_5')
// (7, 13, 'local_g1_5')
// (7, 13, 'lutff_0/in_3')
// (7, 13, 'lutff_1/in_2')
// (7, 13, 'lutff_6/in_2')
// (7, 13, 'sp4_h_r_21')
// (7, 13, 'sp4_r_v_b_4')
// (7, 14, 'local_g3_1')
// (7, 14, 'lutff_5/in_3')
// (7, 14, 'sp4_r_v_b_41')
// (7, 15, 'sp4_r_v_b_28')
// (7, 16, 'sp4_r_v_b_17')
// (8, 5, 'sp12_h_l_23')
// (8, 5, 'sp12_v_t_23')
// (8, 6, 'sp12_v_b_23')
// (8, 7, 'sp12_v_b_20')
// (8, 7, 'sp4_h_r_26')
// (8, 8, 'sp12_v_b_19')
// (8, 9, 'local_g2_1')
// (8, 9, 'lutff_1/in_2')
// (8, 9, 'lutff_2/in_3')
// (8, 9, 'lutff_7/in_2')
// (8, 9, 'sp12_v_b_16')
// (8, 9, 'sp4_h_l_47')
// (8, 9, 'sp4_h_r_25')
// (8, 9, 'sp4_v_t_41')
// (8, 10, 'local_g3_7')
// (8, 10, 'lutff_1/in_3')
// (8, 10, 'sp12_v_b_15')
// (8, 10, 'sp4_v_b_41')
// (8, 11, 'sp12_v_b_12')
// (8, 11, 'sp4_v_b_28')
// (8, 12, 'local_g3_3')
// (8, 12, 'lutff_0/in_2')
// (8, 12, 'sp12_v_b_11')
// (8, 12, 'sp4_v_b_17')
// (8, 13, 'local_g2_0')
// (8, 13, 'lutff_1/in_3')
// (8, 13, 'lutff_5/in_3')
// (8, 13, 'lutff_6/in_2')
// (8, 13, 'sp12_v_b_8')
// (8, 13, 'sp4_h_r_32')
// (8, 13, 'sp4_v_b_4')
// (8, 13, 'sp4_v_t_41')
// (8, 14, 'sp12_v_b_7')
// (8, 14, 'sp4_v_b_41')
// (8, 15, 'sp12_v_b_4')
// (8, 15, 'sp4_v_b_28')
// (8, 16, 'sp12_v_b_3')
// (8, 16, 'sp4_v_b_17')
// (8, 17, 'span12_vert_0')
// (8, 17, 'span4_vert_4')
// (9, 7, 'sp4_h_r_39')
// (9, 9, 'sp4_h_r_36')
// (9, 13, 'sp4_h_r_45')
// (10, 7, 'sp4_h_l_39')
// (10, 9, 'sp4_h_l_36')
// (10, 13, 'sp4_h_l_45')

reg n19 = 0;
// (0, 5, 'span4_horz_10')
// (1, 4, 'neigh_op_tnr_1')
// (1, 5, 'neigh_op_rgt_1')
// (1, 5, 'sp4_h_r_23')
// (1, 6, 'neigh_op_bnr_1')
// (1, 8, 'local_g3_0')
// (1, 8, 'lutff_0/in_3')
// (1, 8, 'sp4_r_v_b_40')
// (1, 9, 'sp4_r_v_b_29')
// (1, 10, 'sp4_r_v_b_16')
// (1, 11, 'sp4_r_v_b_5')
// (2, 2, 'sp12_v_t_22')
// (2, 3, 'sp12_v_b_22')
// (2, 4, 'neigh_op_top_1')
// (2, 4, 'sp12_v_b_21')
// (2, 5, 'lutff_1/out')
// (2, 5, 'sp12_v_b_18')
// (2, 5, 'sp4_h_r_34')
// (2, 6, 'neigh_op_bot_1')
// (2, 6, 'sp12_v_b_17')
// (2, 7, 'sp12_v_b_14')
// (2, 7, 'sp4_v_t_40')
// (2, 8, 'local_g2_5')
// (2, 8, 'local_g3_5')
// (2, 8, 'lutff_0/in_3')
// (2, 8, 'lutff_3/in_3')
// (2, 8, 'lutff_7/in_3')
// (2, 8, 'sp12_v_b_13')
// (2, 8, 'sp4_v_b_40')
// (2, 9, 'sp12_v_b_10')
// (2, 9, 'sp4_v_b_29')
// (2, 10, 'sp12_v_b_9')
// (2, 10, 'sp4_v_b_16')
// (2, 11, 'sp12_v_b_6')
// (2, 11, 'sp4_h_r_11')
// (2, 11, 'sp4_h_r_7')
// (2, 11, 'sp4_v_b_5')
// (2, 12, 'sp12_v_b_5')
// (2, 13, 'sp12_v_b_2')
// (2, 14, 'sp12_v_b_1')
// (3, 4, 'neigh_op_tnl_1')
// (3, 5, 'neigh_op_lft_1')
// (3, 5, 'sp4_h_r_47')
// (3, 6, 'neigh_op_bnl_1')
// (3, 6, 'sp4_r_v_b_47')
// (3, 7, 'sp4_r_v_b_34')
// (3, 8, 'sp4_r_v_b_23')
// (3, 9, 'sp4_r_v_b_10')
// (3, 10, 'sp4_r_v_b_43')
// (3, 11, 'sp4_h_r_18')
// (3, 11, 'sp4_h_r_22')
// (3, 11, 'sp4_r_v_b_30')
// (3, 12, 'sp4_r_v_b_19')
// (3, 13, 'sp4_r_v_b_6')
// (4, 5, 'sp4_h_l_47')
// (4, 5, 'sp4_v_t_47')
// (4, 6, 'sp4_v_b_47')
// (4, 7, 'sp4_v_b_34')
// (4, 8, 'local_g0_7')
// (4, 8, 'lutff_0/in_3')
// (4, 8, 'sp4_v_b_23')
// (4, 9, 'local_g1_2')
// (4, 9, 'lutff_0/in_3')
// (4, 9, 'lutff_4/in_3')
// (4, 9, 'lutff_6/in_3')
// (4, 9, 'sp4_h_r_11')
// (4, 9, 'sp4_h_r_4')
// (4, 9, 'sp4_v_b_10')
// (4, 9, 'sp4_v_t_43')
// (4, 10, 'local_g2_3')
// (4, 10, 'local_g3_3')
// (4, 10, 'lutff_2/in_3')
// (4, 10, 'lutff_3/in_3')
// (4, 10, 'sp4_v_b_43')
// (4, 11, 'sp4_h_r_31')
// (4, 11, 'sp4_h_r_35')
// (4, 11, 'sp4_v_b_30')
// (4, 12, 'sp4_v_b_19')
// (4, 13, 'sp4_v_b_6')
// (5, 8, 'sp4_r_v_b_42')
// (5, 9, 'sp4_h_r_17')
// (5, 9, 'sp4_h_r_22')
// (5, 9, 'sp4_r_v_b_31')
// (5, 10, 'sp4_r_v_b_18')
// (5, 11, 'local_g1_7')
// (5, 11, 'local_g3_6')
// (5, 11, 'lutff_0/in_3')
// (5, 11, 'lutff_4/in_3')
// (5, 11, 'lutff_7/in_3')
// (5, 11, 'sp4_h_r_42')
// (5, 11, 'sp4_h_r_46')
// (5, 11, 'sp4_r_v_b_7')
// (6, 7, 'sp4_v_t_42')
// (6, 8, 'sp4_v_b_42')
// (6, 9, 'local_g2_4')
// (6, 9, 'local_g3_4')
// (6, 9, 'lutff_1/in_3')
// (6, 9, 'lutff_2/in_3')
// (6, 9, 'lutff_4/in_3')
// (6, 9, 'sp4_h_r_28')
// (6, 9, 'sp4_h_r_35')
// (6, 9, 'sp4_v_b_31')
// (6, 10, 'local_g0_2')
// (6, 10, 'local_g1_2')
// (6, 10, 'lutff_0/in_3')
// (6, 10, 'lutff_5/in_3')
// (6, 10, 'lutff_6/in_3')
// (6, 10, 'sp4_v_b_18')
// (6, 11, 'local_g0_3')
// (6, 11, 'local_g1_7')
// (6, 11, 'lutff_0/in_3')
// (6, 11, 'lutff_3/in_3')
// (6, 11, 'lutff_7/in_3')
// (6, 11, 'sp4_h_l_42')
// (6, 11, 'sp4_h_l_46')
// (6, 11, 'sp4_h_r_11')
// (6, 11, 'sp4_v_b_7')
// (7, 6, 'sp4_r_v_b_41')
// (7, 6, 'sp4_r_v_b_46')
// (7, 7, 'sp4_r_v_b_28')
// (7, 7, 'sp4_r_v_b_35')
// (7, 8, 'local_g3_1')
// (7, 8, 'local_g3_6')
// (7, 8, 'lutff_1/in_3')
// (7, 8, 'lutff_4/in_3')
// (7, 8, 'sp4_r_v_b_17')
// (7, 8, 'sp4_r_v_b_22')
// (7, 9, 'local_g2_1')
// (7, 9, 'lutff_0/in_3')
// (7, 9, 'sp4_h_r_41')
// (7, 9, 'sp4_h_r_46')
// (7, 9, 'sp4_r_v_b_11')
// (7, 9, 'sp4_r_v_b_4')
// (7, 11, 'sp4_h_r_22')
// (8, 5, 'sp4_v_t_41')
// (8, 5, 'sp4_v_t_46')
// (8, 6, 'sp4_v_b_41')
// (8, 6, 'sp4_v_b_46')
// (8, 7, 'sp4_v_b_28')
// (8, 7, 'sp4_v_b_35')
// (8, 8, 'sp4_v_b_17')
// (8, 8, 'sp4_v_b_22')
// (8, 9, 'sp4_h_l_41')
// (8, 9, 'sp4_h_l_46')
// (8, 9, 'sp4_v_b_11')
// (8, 9, 'sp4_v_b_4')
// (8, 11, 'sp4_h_r_35')
// (9, 11, 'sp4_h_r_46')
// (10, 11, 'sp4_h_l_46')

reg n20 = 0;
// (0, 6, 'span12_horz_0')
// (1, 5, 'neigh_op_tnr_6')
// (1, 6, 'neigh_op_rgt_6')
// (1, 6, 'sp12_h_r_3')
// (1, 7, 'neigh_op_bnr_6')
// (2, 5, 'neigh_op_top_6')
// (2, 6, 'lutff_6/out')
// (2, 6, 'sp12_h_r_4')
// (2, 7, 'neigh_op_bot_6')
// (3, 5, 'neigh_op_tnl_6')
// (3, 6, 'neigh_op_lft_6')
// (3, 6, 'sp12_h_r_7')
// (3, 7, 'neigh_op_bnl_6')
// (4, 6, 'local_g1_0')
// (4, 6, 'lutff_3/in_0')
// (4, 6, 'sp12_h_r_8')
// (5, 6, 'sp12_h_r_11')
// (6, 6, 'sp12_h_r_12')
// (7, 6, 'sp12_h_r_15')
// (8, 6, 'sp12_h_r_16')
// (9, 6, 'sp12_h_r_19')
// (10, 6, 'sp12_h_r_20')
// (11, 6, 'sp12_h_r_23')
// (12, 6, 'sp12_h_l_23')

reg n21 = 0;
// (0, 6, 'span12_horz_10')
// (1, 5, 'neigh_op_tnr_3')
// (1, 6, 'neigh_op_rgt_3')
// (1, 6, 'sp12_h_r_13')
// (1, 7, 'neigh_op_bnr_3')
// (2, 5, 'neigh_op_top_3')
// (2, 6, 'lutff_3/out')
// (2, 6, 'sp12_h_r_14')
// (2, 7, 'neigh_op_bot_3')
// (3, 5, 'neigh_op_tnl_3')
// (3, 6, 'neigh_op_lft_3')
// (3, 6, 'sp12_h_r_17')
// (3, 7, 'neigh_op_bnl_3')
// (4, 6, 'local_g0_2')
// (4, 6, 'lutff_4/in_0')
// (4, 6, 'sp12_h_r_18')
// (5, 6, 'sp12_h_r_21')
// (6, 6, 'sp12_h_r_22')
// (7, 6, 'sp12_h_l_22')

wire n22;
// (0, 6, 'span12_horz_11')
// (1, 6, 'sp12_h_r_12')
// (2, 6, 'sp12_h_r_15')
// (3, 6, 'sp12_h_r_16')
// (4, 5, 'neigh_op_tnr_6')
// (4, 6, 'neigh_op_rgt_6')
// (4, 6, 'sp12_h_r_19')
// (4, 6, 'sp4_r_v_b_44')
// (4, 7, 'neigh_op_bnr_6')
// (4, 7, 'sp4_r_v_b_33')
// (4, 8, 'sp4_r_v_b_20')
// (4, 9, 'sp4_r_v_b_9')
// (4, 10, 'sp4_r_v_b_44')
// (4, 11, 'sp4_r_v_b_33')
// (4, 12, 'sp4_r_v_b_20')
// (4, 13, 'sp4_r_v_b_9')
// (5, 5, 'neigh_op_top_6')
// (5, 5, 'sp4_v_t_44')
// (5, 6, 'lutff_6/out')
// (5, 6, 'sp12_h_r_20')
// (5, 6, 'sp4_v_b_44')
// (5, 7, 'neigh_op_bot_6')
// (5, 7, 'sp4_v_b_33')
// (5, 8, 'sp4_v_b_20')
// (5, 9, 'local_g0_1')
// (5, 9, 'lutff_1/in_2')
// (5, 9, 'sp4_v_b_9')
// (5, 9, 'sp4_v_t_44')
// (5, 10, 'sp4_v_b_44')
// (5, 11, 'local_g2_1')
// (5, 11, 'lutff_2/in_3')
// (5, 11, 'lutff_6/in_3')
// (5, 11, 'sp4_v_b_33')
// (5, 12, 'sp4_v_b_20')
// (5, 13, 'sp4_v_b_9')
// (6, 5, 'neigh_op_tnl_6')
// (6, 6, 'neigh_op_lft_6')
// (6, 6, 'sp12_h_r_23')
// (6, 7, 'neigh_op_bnl_6')
// (7, 6, 'sp12_h_l_23')
// (7, 6, 'sp12_v_t_23')
// (7, 7, 'sp12_v_b_23')
// (7, 8, 'sp12_v_b_20')
// (7, 9, 'sp12_v_b_19')
// (7, 10, 'sp12_v_b_16')
// (7, 11, 'local_g3_7')
// (7, 11, 'lutff_7/in_3')
// (7, 11, 'sp12_v_b_15')
// (7, 12, 'sp12_v_b_12')
// (7, 13, 'sp12_v_b_11')
// (7, 14, 'sp12_v_b_8')
// (7, 15, 'sp12_v_b_7')
// (7, 16, 'sp12_v_b_4')
// (7, 17, 'span12_vert_3')

wire n23;
// (0, 6, 'span12_horz_13')
// (1, 6, 'sp12_h_r_14')
// (2, 6, 'sp12_h_r_17')
// (3, 6, 'sp12_h_r_18')
// (4, 5, 'neigh_op_tnr_7')
// (4, 6, 'neigh_op_rgt_7')
// (4, 6, 'sp12_h_r_21')
// (4, 7, 'neigh_op_bnr_7')
// (5, 5, 'neigh_op_top_7')
// (5, 6, 'local_g1_6')
// (5, 6, 'lutff_6/in_3')
// (5, 6, 'lutff_7/out')
// (5, 6, 'sp12_h_r_22')
// (5, 7, 'local_g0_7')
// (5, 7, 'local_g1_7')
// (5, 7, 'lutff_0/in_3')
// (5, 7, 'lutff_1/in_3')
// (5, 7, 'neigh_op_bot_7')
// (6, 5, 'neigh_op_tnl_7')
// (6, 6, 'neigh_op_lft_7')
// (6, 6, 'sp12_h_l_22')
// (6, 7, 'neigh_op_bnl_7')

reg n24 = 0;
// (0, 6, 'span12_horz_2')
// (1, 6, 'sp12_h_r_5')
// (2, 6, 'sp12_h_r_6')
// (3, 5, 'neigh_op_tnr_1')
// (3, 6, 'neigh_op_rgt_1')
// (3, 6, 'sp12_h_r_9')
// (3, 7, 'neigh_op_bnr_1')
// (4, 3, 'sp12_v_t_22')
// (4, 4, 'sp12_v_b_22')
// (4, 5, 'neigh_op_top_1')
// (4, 5, 'sp12_v_b_21')
// (4, 6, 'lutff_1/out')
// (4, 6, 'sp12_h_r_10')
// (4, 6, 'sp12_v_b_18')
// (4, 6, 'sp4_h_r_2')
// (4, 7, 'neigh_op_bot_1')
// (4, 7, 'sp12_v_b_17')
// (4, 8, 'sp12_v_b_14')
// (4, 9, 'sp12_v_b_13')
// (4, 10, 'local_g3_2')
// (4, 10, 'lutff_7/in_2')
// (4, 10, 'sp12_v_b_10')
// (4, 11, 'local_g2_1')
// (4, 11, 'lutff_3/in_2')
// (4, 11, 'sp12_v_b_9')
// (4, 12, 'sp12_v_b_6')
// (4, 13, 'sp12_v_b_5')
// (4, 14, 'sp12_v_b_2')
// (4, 15, 'sp12_v_b_1')
// (5, 5, 'neigh_op_tnl_1')
// (5, 6, 'neigh_op_lft_1')
// (5, 6, 'sp12_h_r_13')
// (5, 6, 'sp4_h_r_15')
// (5, 7, 'neigh_op_bnl_1')
// (6, 6, 'sp12_h_r_14')
// (6, 6, 'sp4_h_r_26')
// (7, 6, 'sp12_h_r_17')
// (7, 6, 'sp4_h_r_39')
// (7, 7, 'sp4_r_v_b_39')
// (7, 8, 'sp4_r_v_b_26')
// (7, 9, 'sp4_r_v_b_15')
// (7, 10, 'sp4_r_v_b_2')
// (7, 11, 'sp4_r_v_b_39')
// (7, 12, 'sp4_r_v_b_26')
// (7, 13, 'sp4_r_v_b_15')
// (7, 14, 'sp4_r_v_b_2')
// (8, 6, 'local_g0_2')
// (8, 6, 'lutff_6/in_0')
// (8, 6, 'sp12_h_r_18')
// (8, 6, 'sp4_h_l_39')
// (8, 6, 'sp4_v_t_39')
// (8, 7, 'sp4_v_b_39')
// (8, 8, 'sp4_v_b_26')
// (8, 9, 'sp4_v_b_15')
// (8, 10, 'sp4_v_b_2')
// (8, 10, 'sp4_v_t_39')
// (8, 11, 'sp4_v_b_39')
// (8, 12, 'sp4_v_b_26')
// (8, 13, 'local_g0_7')
// (8, 13, 'lutff_7/in_0')
// (8, 13, 'sp4_v_b_15')
// (8, 14, 'sp4_v_b_2')
// (9, 6, 'sp12_h_r_21')
// (10, 6, 'sp12_h_r_22')
// (11, 6, 'sp12_h_l_22')

wire n25;
// (0, 6, 'span4_horz_11')
// (1, 6, 'sp4_h_r_22')
// (2, 6, 'local_g2_3')
// (2, 6, 'lutff_3/in_0')
// (2, 6, 'sp4_h_r_35')
// (3, 2, 'neigh_op_tnr_7')
// (3, 2, 'sp4_r_v_b_43')
// (3, 3, 'neigh_op_rgt_7')
// (3, 3, 'sp4_r_v_b_30')
// (3, 3, 'sp4_r_v_b_46')
// (3, 4, 'neigh_op_bnr_7')
// (3, 4, 'sp4_r_v_b_19')
// (3, 4, 'sp4_r_v_b_35')
// (3, 5, 'sp4_r_v_b_22')
// (3, 5, 'sp4_r_v_b_6')
// (3, 6, 'sp4_h_r_46')
// (3, 6, 'sp4_r_v_b_11')
// (4, 1, 'sp4_v_t_43')
// (4, 2, 'neigh_op_top_7')
// (4, 2, 'sp4_v_b_43')
// (4, 2, 'sp4_v_t_46')
// (4, 3, 'lutff_7/out')
// (4, 3, 'sp4_v_b_30')
// (4, 3, 'sp4_v_b_46')
// (4, 4, 'neigh_op_bot_7')
// (4, 4, 'sp4_v_b_19')
// (4, 4, 'sp4_v_b_35')
// (4, 5, 'local_g1_6')
// (4, 5, 'lutff_7/in_2')
// (4, 5, 'sp4_v_b_22')
// (4, 5, 'sp4_v_b_6')
// (4, 6, 'local_g1_3')
// (4, 6, 'lutff_0/in_2')
// (4, 6, 'sp4_h_l_46')
// (4, 6, 'sp4_v_b_11')
// (5, 2, 'neigh_op_tnl_7')
// (5, 3, 'neigh_op_lft_7')
// (5, 4, 'neigh_op_bnl_7')

reg n26 = 0;
// (0, 7, 'logic_op_tnr_2')
// (0, 8, 'logic_op_rgt_2')
// (0, 9, 'logic_op_bnr_2')
// (1, 5, 'sp4_r_v_b_40')
// (1, 6, 'sp4_r_v_b_29')
// (1, 7, 'neigh_op_top_2')
// (1, 7, 'sp4_r_v_b_16')
// (1, 8, 'lutff_2/out')
// (1, 8, 'sp4_r_v_b_5')
// (1, 9, 'neigh_op_bot_2')
// (2, 4, 'sp4_v_t_40')
// (2, 5, 'sp4_v_b_40')
// (2, 6, 'sp4_v_b_29')
// (2, 7, 'neigh_op_tnl_2')
// (2, 7, 'sp4_v_b_16')
// (2, 8, 'local_g1_5')
// (2, 8, 'lutff_7/in_1')
// (2, 8, 'neigh_op_lft_2')
// (2, 8, 'sp4_v_b_5')
// (2, 9, 'neigh_op_bnl_2')

reg n27 = 0;
// (0, 7, 'span12_horz_10')
// (1, 6, 'neigh_op_tnr_3')
// (1, 7, 'neigh_op_rgt_3')
// (1, 7, 'sp12_h_r_13')
// (1, 8, 'neigh_op_bnr_3')
// (2, 6, 'neigh_op_top_3')
// (2, 7, 'lutff_3/out')
// (2, 7, 'sp12_h_r_14')
// (2, 8, 'neigh_op_bot_3')
// (3, 6, 'neigh_op_tnl_3')
// (3, 7, 'neigh_op_lft_3')
// (3, 7, 'sp12_h_r_17')
// (3, 8, 'neigh_op_bnl_3')
// (4, 7, 'local_g0_2')
// (4, 7, 'lutff_4/in_0')
// (4, 7, 'sp12_h_r_18')
// (5, 7, 'sp12_h_r_21')
// (6, 7, 'sp12_h_r_22')
// (7, 7, 'sp12_h_l_22')

reg n28 = 0;
// (0, 7, 'span12_horz_7')
// (1, 7, 'sp12_h_r_8')
// (2, 7, 'local_g0_3')
// (2, 7, 'lutff_3/in_0')
// (2, 7, 'sp12_h_r_11')
// (3, 7, 'sp12_h_r_12')
// (4, 6, 'neigh_op_tnr_4')
// (4, 7, 'neigh_op_rgt_4')
// (4, 7, 'sp12_h_r_15')
// (4, 8, 'neigh_op_bnr_4')
// (5, 6, 'neigh_op_top_4')
// (5, 7, 'lutff_4/out')
// (5, 7, 'sp12_h_r_16')
// (5, 8, 'neigh_op_bot_4')
// (6, 6, 'neigh_op_tnl_4')
// (6, 7, 'neigh_op_lft_4')
// (6, 7, 'sp12_h_r_19')
// (6, 8, 'neigh_op_bnl_4')
// (7, 7, 'sp12_h_r_20')
// (8, 7, 'sp12_h_r_23')
// (9, 7, 'sp12_h_l_23')

reg n29 = 0;
// (0, 7, 'span12_horz_9')
// (1, 7, 'sp12_h_r_10')
// (2, 7, 'sp12_h_r_13')
// (3, 7, 'sp12_h_r_14')
// (4, 7, 'sp12_h_r_17')
// (5, 7, 'sp12_h_r_18')
// (5, 7, 'sp4_h_r_6')
// (6, 6, 'neigh_op_tnr_7')
// (6, 7, 'local_g0_5')
// (6, 7, 'local_g1_3')
// (6, 7, 'lutff_2/in_2')
// (6, 7, 'lutff_7/in_2')
// (6, 7, 'neigh_op_rgt_7')
// (6, 7, 'sp12_h_r_21')
// (6, 7, 'sp4_h_r_19')
// (6, 8, 'neigh_op_bnr_7')
// (7, 6, 'neigh_op_top_7')
// (7, 7, 'lutff_7/out')
// (7, 7, 'sp12_h_r_22')
// (7, 7, 'sp4_h_r_30')
// (7, 8, 'neigh_op_bot_7')
// (8, 6, 'neigh_op_tnl_7')
// (8, 7, 'local_g1_7')
// (8, 7, 'lutff_6/in_0')
// (8, 7, 'neigh_op_lft_7')
// (8, 7, 'sp12_h_l_22')
// (8, 7, 'sp4_h_r_43')
// (8, 8, 'neigh_op_bnl_7')
// (8, 8, 'sp4_r_v_b_46')
// (8, 9, 'sp4_r_v_b_35')
// (8, 10, 'sp4_r_v_b_22')
// (8, 11, 'sp4_r_v_b_11')
// (9, 7, 'sp4_h_l_43')
// (9, 7, 'sp4_v_t_46')
// (9, 8, 'local_g2_6')
// (9, 8, 'lutff_6/in_0')
// (9, 8, 'sp4_v_b_46')
// (9, 9, 'sp4_v_b_35')
// (9, 10, 'sp4_v_b_22')
// (9, 11, 'sp4_v_b_11')

wire n30;
// (0, 8, 'span12_horz_0')
// (1, 8, 'sp12_h_r_3')
// (2, 8, 'sp12_h_r_4')
// (3, 7, 'neigh_op_tnr_0')
// (3, 8, 'neigh_op_rgt_0')
// (3, 8, 'sp12_h_r_7')
// (3, 9, 'neigh_op_bnr_0')
// (4, 7, 'neigh_op_top_0')
// (4, 8, 'lutff_0/out')
// (4, 8, 'sp12_h_r_8')
// (4, 9, 'neigh_op_bot_0')
// (5, 7, 'neigh_op_tnl_0')
// (5, 8, 'neigh_op_lft_0')
// (5, 8, 'sp12_h_r_11')
// (5, 9, 'neigh_op_bnl_0')
// (6, 8, 'local_g0_4')
// (6, 8, 'lutff_3/in_1')
// (6, 8, 'sp12_h_r_12')
// (7, 8, 'local_g1_7')
// (7, 8, 'lutff_7/in_1')
// (7, 8, 'sp12_h_r_15')
// (8, 8, 'sp12_h_r_16')
// (9, 8, 'sp12_h_r_19')
// (10, 8, 'sp12_h_r_20')
// (11, 8, 'sp12_h_r_23')
// (12, 8, 'sp12_h_l_23')

reg n31 = 0;
// (0, 8, 'span12_horz_2')
// (1, 8, 'local_g1_5')
// (1, 8, 'lutff_2/in_0')
// (1, 8, 'sp12_h_r_5')
// (2, 8, 'sp12_h_r_6')
// (3, 7, 'neigh_op_tnr_1')
// (3, 8, 'neigh_op_rgt_1')
// (3, 8, 'sp12_h_r_9')
// (3, 9, 'neigh_op_bnr_1')
// (4, 7, 'neigh_op_top_1')
// (4, 8, 'local_g0_1')
// (4, 8, 'lutff_1/out')
// (4, 8, 'lutff_6/in_1')
// (4, 8, 'sp12_h_r_10')
// (4, 9, 'neigh_op_bot_1')
// (5, 7, 'neigh_op_tnl_1')
// (5, 8, 'neigh_op_lft_1')
// (5, 8, 'sp12_h_r_13')
// (5, 9, 'neigh_op_bnl_1')
// (6, 8, 'sp12_h_r_14')
// (7, 8, 'sp12_h_r_17')
// (8, 8, 'sp12_h_r_18')
// (9, 8, 'sp12_h_r_21')
// (10, 8, 'sp12_h_r_22')
// (11, 8, 'sp12_h_l_22')

wire n32;
// (0, 8, 'span12_horz_3')
// (1, 8, 'sp12_h_r_4')
// (2, 8, 'sp12_h_r_7')
// (3, 8, 'sp12_h_r_8')
// (4, 7, 'neigh_op_tnr_2')
// (4, 8, 'neigh_op_rgt_2')
// (4, 8, 'sp12_h_r_11')
// (4, 9, 'neigh_op_bnr_2')
// (5, 7, 'neigh_op_top_2')
// (5, 8, 'lutff_2/out')
// (5, 8, 'sp12_h_r_12')
// (5, 9, 'neigh_op_bot_2')
// (6, 7, 'neigh_op_tnl_2')
// (6, 8, 'neigh_op_lft_2')
// (6, 8, 'sp12_h_r_15')
// (6, 8, 'sp4_h_r_9')
// (6, 9, 'neigh_op_bnl_2')
// (7, 8, 'local_g0_4')
// (7, 8, 'local_g1_0')
// (7, 8, 'lutff_0/in_3')
// (7, 8, 'lutff_2/in_3')
// (7, 8, 'lutff_5/in_3')
// (7, 8, 'sp12_h_r_16')
// (7, 8, 'sp4_h_r_20')
// (8, 8, 'sp12_h_r_19')
// (8, 8, 'sp4_h_r_33')
// (9, 8, 'local_g0_4')
// (9, 8, 'lutff_3/in_3')
// (9, 8, 'sp12_h_r_20')
// (9, 8, 'sp4_h_r_44')
// (10, 8, 'sp12_h_r_23')
// (10, 8, 'sp4_h_l_44')
// (11, 8, 'sp12_h_l_23')

reg n33 = 0;
// (0, 8, 'span12_horz_4')
// (1, 8, 'sp12_h_r_7')
// (2, 8, 'local_g1_0')
// (2, 8, 'lutff_3/in_2')
// (2, 8, 'sp12_h_r_8')
// (3, 7, 'neigh_op_tnr_2')
// (3, 8, 'neigh_op_rgt_2')
// (3, 8, 'sp12_h_r_11')
// (3, 9, 'neigh_op_bnr_2')
// (4, 7, 'neigh_op_top_2')
// (4, 8, 'local_g1_2')
// (4, 8, 'lutff_2/out')
// (4, 8, 'lutff_4/in_1')
// (4, 8, 'sp12_h_r_12')
// (4, 9, 'neigh_op_bot_2')
// (5, 7, 'neigh_op_tnl_2')
// (5, 8, 'neigh_op_lft_2')
// (5, 8, 'sp12_h_r_15')
// (5, 9, 'neigh_op_bnl_2')
// (6, 8, 'sp12_h_r_16')
// (7, 8, 'sp12_h_r_19')
// (8, 8, 'sp12_h_r_20')
// (9, 8, 'sp12_h_r_23')
// (10, 8, 'sp12_h_l_23')

reg n34 = 0;
// (0, 8, 'span4_horz_8')
// (1, 7, 'neigh_op_tnr_0')
// (1, 8, 'neigh_op_rgt_0')
// (1, 8, 'sp4_h_r_21')
// (1, 9, 'neigh_op_bnr_0')
// (2, 7, 'neigh_op_top_0')
// (2, 8, 'lutff_0/out')
// (2, 8, 'sp4_h_r_32')
// (2, 9, 'neigh_op_bot_0')
// (3, 5, 'sp4_r_v_b_45')
// (3, 6, 'sp4_r_v_b_32')
// (3, 7, 'neigh_op_tnl_0')
// (3, 7, 'sp4_r_v_b_21')
// (3, 8, 'neigh_op_lft_0')
// (3, 8, 'sp4_h_r_45')
// (3, 8, 'sp4_r_v_b_8')
// (3, 9, 'neigh_op_bnl_0')
// (4, 4, 'sp4_v_t_45')
// (4, 5, 'sp4_v_b_45')
// (4, 6, 'sp4_v_b_32')
// (4, 7, 'sp4_v_b_21')
// (4, 8, 'local_g1_0')
// (4, 8, 'lutff_0/in_1')
// (4, 8, 'sp4_h_l_45')
// (4, 8, 'sp4_v_b_8')

reg n35 = 0;
// (0, 9, 'logic_op_tnr_5')
// (0, 10, 'logic_op_rgt_5')
// (0, 11, 'logic_op_bnr_5')
// (1, 9, 'neigh_op_top_5')
// (1, 10, 'lutff_5/out')
// (1, 11, 'neigh_op_bot_5')
// (2, 9, 'neigh_op_tnl_5')
// (2, 10, 'local_g0_5')
// (2, 10, 'lutff_1/in_0')
// (2, 10, 'neigh_op_lft_5')
// (2, 11, 'neigh_op_bnl_5')

reg n36 = 0;
// (0, 9, 'span12_horz_14')
// (1, 9, 'sp12_h_r_17')
// (2, 9, 'local_g1_2')
// (2, 9, 'lutff_5/in_0')
// (2, 9, 'sp12_h_r_18')
// (3, 8, 'neigh_op_tnr_7')
// (3, 9, 'neigh_op_rgt_7')
// (3, 9, 'sp12_h_r_21')
// (3, 10, 'neigh_op_bnr_7')
// (4, 8, 'neigh_op_top_7')
// (4, 9, 'local_g0_7')
// (4, 9, 'lutff_2/in_1')
// (4, 9, 'lutff_7/out')
// (4, 9, 'sp12_h_r_22')
// (4, 10, 'neigh_op_bot_7')
// (5, 8, 'neigh_op_tnl_7')
// (5, 9, 'neigh_op_lft_7')
// (5, 9, 'sp12_h_l_22')
// (5, 10, 'neigh_op_bnl_7')

reg n37 = 0;
// (0, 9, 'span12_horz_5')
// (1, 9, 'sp12_h_r_6')
// (2, 9, 'sp12_h_r_9')
// (3, 9, 'sp12_h_r_10')
// (4, 9, 'sp12_h_r_13')
// (5, 9, 'local_g1_6')
// (5, 9, 'lutff_5/in_0')
// (5, 9, 'sp12_h_r_14')
// (6, 8, 'neigh_op_tnr_5')
// (6, 9, 'neigh_op_rgt_5')
// (6, 9, 'sp12_h_r_17')
// (6, 10, 'neigh_op_bnr_5')
// (7, 8, 'neigh_op_top_5')
// (7, 9, 'lutff_5/out')
// (7, 9, 'sp12_h_r_18')
// (7, 10, 'neigh_op_bot_5')
// (8, 8, 'neigh_op_tnl_5')
// (8, 9, 'neigh_op_lft_5')
// (8, 9, 'sp12_h_r_21')
// (8, 10, 'neigh_op_bnl_5')
// (9, 9, 'sp12_h_r_22')
// (10, 9, 'sp12_h_l_22')

reg n38 = 0;
// (0, 9, 'span12_horz_6')
// (1, 9, 'sp12_h_r_9')
// (2, 9, 'sp12_h_r_10')
// (3, 9, 'sp12_h_r_13')
// (4, 9, 'sp12_h_r_14')
// (5, 9, 'sp12_h_r_17')
// (6, 9, 'sp12_h_r_18')
// (7, 9, 'sp12_h_r_21')
// (7, 9, 'sp4_h_r_10')
// (8, 5, 'neigh_op_tnr_3')
// (8, 6, 'local_g2_3')
// (8, 6, 'lutff_7/in_0')
// (8, 6, 'neigh_op_rgt_3')
// (8, 7, 'neigh_op_bnr_3')
// (8, 9, 'local_g0_6')
// (8, 9, 'local_g0_7')
// (8, 9, 'lutff_0/in_2')
// (8, 9, 'lutff_3/in_2')
// (8, 9, 'sp12_h_r_22')
// (8, 9, 'sp4_h_r_23')
// (9, 0, 'span12_vert_17')
// (9, 1, 'sp12_v_b_17')
// (9, 2, 'sp12_v_b_14')
// (9, 3, 'sp12_v_b_13')
// (9, 4, 'sp12_v_b_10')
// (9, 5, 'neigh_op_top_3')
// (9, 5, 'sp12_v_b_9')
// (9, 6, 'lutff_3/out')
// (9, 6, 'sp12_v_b_6')
// (9, 7, 'neigh_op_bot_3')
// (9, 7, 'sp12_v_b_5')
// (9, 8, 'sp12_v_b_2')
// (9, 9, 'local_g3_2')
// (9, 9, 'lutff_5/in_0')
// (9, 9, 'sp12_h_l_22')
// (9, 9, 'sp12_v_b_1')
// (9, 9, 'sp4_h_r_34')
// (10, 5, 'neigh_op_tnl_3')
// (10, 6, 'neigh_op_lft_3')
// (10, 7, 'neigh_op_bnl_3')
// (10, 9, 'sp4_h_r_47')
// (11, 9, 'sp4_h_l_47')

wire n39;
// (0, 10, 'span12_horz_0')
// (1, 10, 'sp12_h_r_3')
// (2, 10, 'sp12_h_r_4')
// (3, 8, 'sp4_r_v_b_40')
// (3, 9, 'neigh_op_tnr_0')
// (3, 9, 'sp4_r_v_b_29')
// (3, 10, 'neigh_op_rgt_0')
// (3, 10, 'sp12_h_r_7')
// (3, 10, 'sp4_r_v_b_16')
// (3, 11, 'neigh_op_bnr_0')
// (3, 11, 'sp4_r_v_b_5')
// (4, 7, 'sp4_v_t_40')
// (4, 8, 'sp4_r_v_b_41')
// (4, 8, 'sp4_v_b_40')
// (4, 9, 'neigh_op_top_0')
// (4, 9, 'sp4_r_v_b_28')
// (4, 9, 'sp4_r_v_b_44')
// (4, 9, 'sp4_v_b_29')
// (4, 10, 'local_g1_0')
// (4, 10, 'lutff_0/out')
// (4, 10, 'lutff_7/in_0')
// (4, 10, 'sp12_h_r_8')
// (4, 10, 'sp4_r_v_b_17')
// (4, 10, 'sp4_r_v_b_33')
// (4, 10, 'sp4_v_b_16')
// (4, 11, 'local_g1_5')
// (4, 11, 'lutff_3/in_3')
// (4, 11, 'neigh_op_bot_0')
// (4, 11, 'sp4_h_r_5')
// (4, 11, 'sp4_r_v_b_20')
// (4, 11, 'sp4_r_v_b_4')
// (4, 11, 'sp4_v_b_5')
// (4, 12, 'sp4_r_v_b_9')
// (5, 7, 'sp4_h_r_9')
// (5, 7, 'sp4_v_t_41')
// (5, 8, 'sp4_h_r_2')
// (5, 8, 'sp4_v_b_41')
// (5, 8, 'sp4_v_t_44')
// (5, 9, 'local_g2_0')
// (5, 9, 'lutff_0/in_0')
// (5, 9, 'neigh_op_tnl_0')
// (5, 9, 'sp4_v_b_28')
// (5, 9, 'sp4_v_b_44')
// (5, 10, 'local_g1_1')
// (5, 10, 'lutff_3/in_3')
// (5, 10, 'neigh_op_lft_0')
// (5, 10, 'sp12_h_r_11')
// (5, 10, 'sp4_v_b_17')
// (5, 10, 'sp4_v_b_33')
// (5, 11, 'neigh_op_bnl_0')
// (5, 11, 'sp4_h_r_16')
// (5, 11, 'sp4_v_b_20')
// (5, 11, 'sp4_v_b_4')
// (5, 12, 'local_g1_1')
// (5, 12, 'lutff_4/in_0')
// (5, 12, 'lutff_5/in_3')
// (5, 12, 'sp4_h_r_9')
// (5, 12, 'sp4_v_b_9')
// (6, 7, 'local_g0_4')
// (6, 7, 'lutff_2/in_0')
// (6, 7, 'lutff_7/in_3')
// (6, 7, 'sp4_h_r_20')
// (6, 8, 'local_g0_7')
// (6, 8, 'lutff_3/in_0')
// (6, 8, 'sp4_h_r_15')
// (6, 10, 'sp12_h_r_12')
// (6, 11, 'sp4_h_r_29')
// (6, 12, 'sp4_h_r_20')
// (7, 7, 'sp4_h_r_33')
// (7, 8, 'local_g2_2')
// (7, 8, 'lutff_7/in_3')
// (7, 8, 'sp4_h_r_26')
// (7, 10, 'local_g1_7')
// (7, 10, 'lutff_0/in_0')
// (7, 10, 'sp12_h_r_15')
// (7, 11, 'local_g2_0')
// (7, 11, 'lutff_2/in_0')
// (7, 11, 'sp4_h_r_40')
// (7, 12, 'local_g2_1')
// (7, 12, 'lutff_4/in_3')
// (7, 12, 'sp4_h_r_33')
// (8, 7, 'sp4_h_r_44')
// (8, 8, 'sp4_h_r_39')
// (8, 8, 'sp4_r_v_b_39')
// (8, 9, 'local_g0_2')
// (8, 9, 'lutff_0/in_0')
// (8, 9, 'lutff_3/in_3')
// (8, 9, 'sp4_r_v_b_26')
// (8, 10, 'sp12_h_r_16')
// (8, 10, 'sp4_r_v_b_15')
// (8, 11, 'local_g1_1')
// (8, 11, 'lutff_3/in_3')
// (8, 11, 'sp4_h_l_40')
// (8, 11, 'sp4_h_r_1')
// (8, 11, 'sp4_r_v_b_2')
// (8, 12, 'sp4_h_r_44')
// (9, 7, 'sp4_h_l_44')
// (9, 7, 'sp4_v_t_39')
// (9, 8, 'sp4_h_l_39')
// (9, 8, 'sp4_v_b_39')
// (9, 9, 'sp4_v_b_26')
// (9, 10, 'sp12_h_r_19')
// (9, 10, 'sp4_v_b_15')
// (9, 11, 'sp4_h_r_12')
// (9, 11, 'sp4_v_b_2')
// (9, 12, 'sp4_h_l_44')
// (10, 10, 'sp12_h_r_20')
// (10, 11, 'sp4_h_r_25')
// (11, 10, 'sp12_h_r_23')
// (11, 11, 'sp4_h_r_36')
// (12, 10, 'sp12_h_l_23')
// (12, 11, 'sp4_h_l_36')

reg n40 = 0;
// (0, 10, 'span12_horz_10')
// (1, 9, 'neigh_op_tnr_3')
// (1, 10, 'neigh_op_rgt_3')
// (1, 10, 'sp12_h_r_13')
// (1, 11, 'neigh_op_bnr_3')
// (2, 9, 'neigh_op_top_3')
// (2, 10, 'lutff_3/out')
// (2, 10, 'sp12_h_r_14')
// (2, 11, 'neigh_op_bot_3')
// (3, 9, 'neigh_op_tnl_3')
// (3, 10, 'neigh_op_lft_3')
// (3, 10, 'sp12_h_r_17')
// (3, 11, 'neigh_op_bnl_3')
// (4, 10, 'sp12_h_r_18')
// (5, 10, 'sp12_h_r_21')
// (6, 10, 'sp12_h_r_22')
// (7, 10, 'local_g0_1')
// (7, 10, 'lutff_5/in_0')
// (7, 10, 'sp12_h_l_22')
// (7, 10, 'sp12_h_r_1')
// (8, 7, 'local_g2_7')
// (8, 7, 'lutff_5/in_2')
// (8, 7, 'sp4_r_v_b_39')
// (8, 8, 'sp4_r_v_b_26')
// (8, 9, 'sp4_r_v_b_15')
// (8, 10, 'sp12_h_r_2')
// (8, 10, 'sp4_r_v_b_2')
// (9, 6, 'sp4_v_t_39')
// (9, 7, 'sp4_v_b_39')
// (9, 8, 'sp4_v_b_26')
// (9, 9, 'sp4_v_b_15')
// (9, 10, 'sp12_h_r_5')
// (9, 10, 'sp4_h_r_2')
// (9, 10, 'sp4_v_b_2')
// (10, 10, 'sp12_h_r_6')
// (10, 10, 'sp4_h_r_15')
// (11, 10, 'sp12_h_r_9')
// (11, 10, 'sp4_h_r_26')
// (12, 10, 'sp12_h_r_10')
// (12, 10, 'sp4_h_r_39')
// (13, 10, 'span12_horz_10')
// (13, 10, 'span4_horz_39')

reg n41 = 0;
// (0, 10, 'span12_horz_2')
// (1, 9, 'neigh_op_tnr_7')
// (1, 10, 'neigh_op_rgt_7')
// (1, 10, 'sp12_h_r_5')
// (1, 11, 'neigh_op_bnr_7')
// (2, 9, 'neigh_op_top_7')
// (2, 10, 'lutff_7/out')
// (2, 10, 'sp12_h_r_6')
// (2, 10, 'sp4_r_v_b_47')
// (2, 11, 'neigh_op_bot_7')
// (2, 11, 'sp4_r_v_b_34')
// (2, 12, 'sp4_r_v_b_23')
// (2, 13, 'sp4_r_v_b_10')
// (3, 9, 'neigh_op_tnl_7')
// (3, 9, 'sp4_h_r_10')
// (3, 9, 'sp4_v_t_47')
// (3, 10, 'neigh_op_lft_7')
// (3, 10, 'sp12_h_r_9')
// (3, 10, 'sp4_h_r_4')
// (3, 10, 'sp4_v_b_47')
// (3, 11, 'neigh_op_bnl_7')
// (3, 11, 'sp4_v_b_34')
// (3, 12, 'sp4_v_b_23')
// (3, 13, 'sp4_v_b_10')
// (4, 9, 'sp4_h_r_23')
// (4, 10, 'sp12_h_r_10')
// (4, 10, 'sp4_h_r_17')
// (5, 9, 'sp4_h_r_34')
// (5, 10, 'sp12_h_r_13')
// (5, 10, 'sp4_h_r_28')
// (6, 9, 'local_g2_7')
// (6, 9, 'lutff_0/in_1')
// (6, 9, 'sp4_h_r_47')
// (6, 10, 'local_g2_1')
// (6, 10, 'lutff_4/in_1')
// (6, 10, 'sp12_h_r_14')
// (6, 10, 'sp4_h_r_41')
// (7, 9, 'sp4_h_l_47')
// (7, 10, 'sp12_h_r_17')
// (7, 10, 'sp4_h_l_41')
// (8, 10, 'sp12_h_r_18')
// (9, 10, 'sp12_h_r_21')
// (10, 10, 'sp12_h_r_22')
// (11, 10, 'sp12_h_l_22')

wire n42;
// (0, 10, 'span12_horz_4')
// (1, 10, 'sp12_h_r_7')
// (2, 10, 'sp12_h_r_8')
// (3, 9, 'neigh_op_tnr_2')
// (3, 10, 'neigh_op_rgt_2')
// (3, 10, 'sp12_h_r_11')
// (3, 11, 'neigh_op_bnr_2')
// (4, 0, 'span12_vert_23')
// (4, 1, 'sp12_v_b_23')
// (4, 2, 'sp12_v_b_20')
// (4, 3, 'sp12_v_b_19')
// (4, 4, 'sp12_v_b_16')
// (4, 5, 'sp12_v_b_15')
// (4, 6, 'sp12_v_b_12')
// (4, 7, 'sp12_v_b_11')
// (4, 8, 'sp12_v_b_8')
// (4, 9, 'neigh_op_top_2')
// (4, 9, 'sp12_v_b_7')
// (4, 10, 'lutff_2/out')
// (4, 10, 'sp12_h_r_12')
// (4, 10, 'sp12_v_b_4')
// (4, 11, 'neigh_op_bot_2')
// (4, 11, 'sp12_v_b_3')
// (4, 12, 'sp12_h_r_0')
// (4, 12, 'sp12_v_b_0')
// (5, 9, 'neigh_op_tnl_2')
// (5, 10, 'neigh_op_lft_2')
// (5, 10, 'sp12_h_r_15')
// (5, 11, 'neigh_op_bnl_2')
// (5, 12, 'sp12_h_r_3')
// (6, 10, 'sp12_h_r_16')
// (6, 12, 'sp12_h_r_4')
// (7, 10, 'local_g0_3')
// (7, 10, 'lutff_0/in_1')
// (7, 10, 'sp12_h_r_19')
// (7, 12, 'local_g0_7')
// (7, 12, 'lutff_4/in_1')
// (7, 12, 'sp12_h_r_7')
// (8, 10, 'sp12_h_r_20')
// (8, 12, 'sp12_h_r_8')
// (9, 10, 'sp12_h_r_23')
// (9, 12, 'sp12_h_r_11')
// (10, 10, 'sp12_h_l_23')
// (10, 12, 'sp12_h_r_12')
// (11, 12, 'sp12_h_r_15')
// (12, 12, 'sp12_h_r_16')
// (13, 12, 'span12_horz_16')

reg n43 = 0;
// (0, 10, 'span12_horz_7')
// (1, 10, 'sp12_h_r_8')
// (2, 10, 'local_g0_3')
// (2, 10, 'lutff_7/in_0')
// (2, 10, 'sp12_h_r_11')
// (3, 10, 'sp12_h_r_12')
// (4, 9, 'neigh_op_tnr_4')
// (4, 10, 'neigh_op_rgt_4')
// (4, 10, 'sp12_h_r_15')
// (4, 11, 'neigh_op_bnr_4')
// (5, 9, 'neigh_op_top_4')
// (5, 10, 'lutff_4/out')
// (5, 10, 'sp12_h_r_16')
// (5, 11, 'neigh_op_bot_4')
// (6, 9, 'neigh_op_tnl_4')
// (6, 10, 'neigh_op_lft_4')
// (6, 10, 'sp12_h_r_19')
// (6, 11, 'neigh_op_bnl_4')
// (7, 10, 'sp12_h_r_20')
// (8, 10, 'sp12_h_r_23')
// (9, 10, 'sp12_h_l_23')

reg d_vld = 0;
// (0, 11, 'logic_op_tnr_5')
// (0, 12, 'logic_op_rgt_5')
// (0, 13, 'logic_op_bnr_5')
// (0, 14, 'io_0/D_OUT_0')
// (0, 14, 'io_0/PAD')
// (0, 14, 'local_g0_0')
// (0, 14, 'span4_horz_32')
// (1, 11, 'neigh_op_top_5')
// (1, 11, 'sp4_r_v_b_38')
// (1, 12, 'lutff_5/out')
// (1, 12, 'sp4_r_v_b_27')
// (1, 13, 'neigh_op_bot_5')
// (1, 13, 'sp4_r_v_b_14')
// (1, 14, 'sp4_h_r_45')
// (1, 14, 'sp4_r_v_b_3')
// (2, 10, 'sp4_v_t_38')
// (2, 11, 'neigh_op_tnl_5')
// (2, 11, 'sp4_v_b_38')
// (2, 12, 'neigh_op_lft_5')
// (2, 12, 'sp4_v_b_27')
// (2, 13, 'neigh_op_bnl_5')
// (2, 13, 'sp4_v_b_14')
// (2, 14, 'sp4_h_l_45')
// (2, 14, 'sp4_v_b_3')

reg n45 = 0;
// (0, 11, 'span12_horz_1')
// (1, 11, 'sp12_h_r_2')
// (2, 11, 'local_g1_5')
// (2, 11, 'lutff_2/in_0')
// (2, 11, 'sp12_h_r_5')
// (3, 11, 'sp12_h_r_6')
// (4, 10, 'neigh_op_tnr_1')
// (4, 11, 'neigh_op_rgt_1')
// (4, 11, 'sp12_h_r_9')
// (4, 12, 'neigh_op_bnr_1')
// (5, 10, 'neigh_op_top_1')
// (5, 11, 'local_g0_1')
// (5, 11, 'lutff_1/out')
// (5, 11, 'lutff_3/in_2')
// (5, 11, 'sp12_h_r_10')
// (5, 12, 'neigh_op_bot_1')
// (6, 10, 'neigh_op_tnl_1')
// (6, 11, 'neigh_op_lft_1')
// (6, 11, 'sp12_h_r_13')
// (6, 12, 'neigh_op_bnl_1')
// (7, 11, 'sp12_h_r_14')
// (8, 11, 'sp12_h_r_17')
// (9, 11, 'sp12_h_r_18')
// (10, 11, 'sp12_h_r_21')
// (11, 11, 'sp12_h_r_22')
// (12, 11, 'sp12_h_l_22')

reg n46 = 0;
// (0, 11, 'span12_horz_17')
// (1, 11, 'sp12_h_r_18')
// (2, 11, 'sp12_h_r_21')
// (2, 11, 'sp4_h_r_10')
// (3, 5, 'neigh_op_tnr_5')
// (3, 5, 'sp4_r_v_b_40')
// (3, 6, 'neigh_op_rgt_5')
// (3, 6, 'sp4_r_v_b_29')
// (3, 7, 'neigh_op_bnr_5')
// (3, 7, 'sp4_r_v_b_16')
// (3, 8, 'sp4_r_v_b_5')
// (3, 11, 'sp12_h_r_22')
// (3, 11, 'sp4_h_r_23')
// (4, 0, 'span12_vert_21')
// (4, 1, 'sp12_v_b_21')
// (4, 2, 'sp12_v_b_18')
// (4, 3, 'sp12_v_b_17')
// (4, 4, 'sp12_v_b_14')
// (4, 4, 'sp4_v_t_40')
// (4, 5, 'neigh_op_top_5')
// (4, 5, 'sp12_v_b_13')
// (4, 5, 'sp4_v_b_40')
// (4, 6, 'lutff_5/out')
// (4, 6, 'sp12_v_b_10')
// (4, 6, 'sp4_v_b_29')
// (4, 7, 'neigh_op_bot_5')
// (4, 7, 'sp12_v_b_9')
// (4, 7, 'sp4_v_b_16')
// (4, 8, 'local_g2_6')
// (4, 8, 'local_g3_6')
// (4, 8, 'lutff_1/in_2')
// (4, 8, 'lutff_2/in_0')
// (4, 8, 'lutff_3/in_2')
// (4, 8, 'lutff_4/in_2')
// (4, 8, 'lutff_5/in_2')
// (4, 8, 'lutff_6/in_0')
// (4, 8, 'lutff_7/in_2')
// (4, 8, 'sp12_v_b_6')
// (4, 8, 'sp4_h_r_5')
// (4, 8, 'sp4_v_b_5')
// (4, 9, 'local_g2_5')
// (4, 9, 'local_g3_5')
// (4, 9, 'lutff_1/in_2')
// (4, 9, 'lutff_2/in_0')
// (4, 9, 'lutff_3/in_2')
// (4, 9, 'lutff_5/in_2')
// (4, 9, 'lutff_7/in_1')
// (4, 9, 'sp12_v_b_5')
// (4, 10, 'sp12_v_b_2')
// (4, 11, 'sp12_h_l_22')
// (4, 11, 'sp12_v_b_1')
// (4, 11, 'sp4_h_r_34')
// (5, 5, 'neigh_op_tnl_5')
// (5, 6, 'neigh_op_lft_5')
// (5, 7, 'neigh_op_bnl_5')
// (5, 8, 'sp4_h_r_16')
// (5, 8, 'sp4_r_v_b_41')
// (5, 8, 'sp4_r_v_b_46')
// (5, 8, 'sp4_r_v_b_47')
// (5, 9, 'sp4_r_v_b_28')
// (5, 9, 'sp4_r_v_b_34')
// (5, 9, 'sp4_r_v_b_35')
// (5, 10, 'sp4_r_v_b_17')
// (5, 10, 'sp4_r_v_b_22')
// (5, 10, 'sp4_r_v_b_23')
// (5, 11, 'local_g2_2')
// (5, 11, 'local_g2_7')
// (5, 11, 'lutff_1/in_2')
// (5, 11, 'lutff_2/in_2')
// (5, 11, 'lutff_3/in_1')
// (5, 11, 'lutff_6/in_2')
// (5, 11, 'sp4_h_r_47')
// (5, 11, 'sp4_r_v_b_10')
// (5, 11, 'sp4_r_v_b_11')
// (5, 11, 'sp4_r_v_b_4')
// (5, 12, 'sp4_r_v_b_38')
// (5, 13, 'sp4_r_v_b_27')
// (5, 14, 'sp4_r_v_b_14')
// (5, 15, 'sp4_r_v_b_3')
// (6, 7, 'sp4_v_t_41')
// (6, 7, 'sp4_v_t_46')
// (6, 7, 'sp4_v_t_47')
// (6, 8, 'sp4_h_r_29')
// (6, 8, 'sp4_v_b_41')
// (6, 8, 'sp4_v_b_46')
// (6, 8, 'sp4_v_b_47')
// (6, 9, 'local_g2_2')
// (6, 9, 'local_g3_2')
// (6, 9, 'lutff_3/in_2')
// (6, 9, 'lutff_5/in_0')
// (6, 9, 'lutff_6/in_2')
// (6, 9, 'lutff_7/in_2')
// (6, 9, 'sp4_v_b_28')
// (6, 9, 'sp4_v_b_34')
// (6, 9, 'sp4_v_b_35')
// (6, 10, 'local_g0_6')
// (6, 10, 'local_g0_7')
// (6, 10, 'lutff_1/in_0')
// (6, 10, 'lutff_2/in_2')
// (6, 10, 'lutff_3/in_2')
// (6, 10, 'lutff_7/in_2')
// (6, 10, 'sp4_v_b_17')
// (6, 10, 'sp4_v_b_22')
// (6, 10, 'sp4_v_b_23')
// (6, 11, 'local_g0_2')
// (6, 11, 'local_g1_4')
// (6, 11, 'lutff_1/in_2')
// (6, 11, 'lutff_2/in_2')
// (6, 11, 'lutff_4/in_2')
// (6, 11, 'lutff_5/in_0')
// (6, 11, 'sp4_h_l_47')
// (6, 11, 'sp4_v_b_10')
// (6, 11, 'sp4_v_b_11')
// (6, 11, 'sp4_v_b_4')
// (6, 11, 'sp4_v_t_38')
// (6, 12, 'sp4_v_b_38')
// (6, 13, 'sp4_v_b_27')
// (6, 14, 'sp4_v_b_14')
// (6, 15, 'sp4_v_b_3')
// (7, 5, 'sp4_r_v_b_46')
// (7, 6, 'sp4_r_v_b_35')
// (7, 7, 'sp4_r_v_b_22')
// (7, 8, 'local_g2_0')
// (7, 8, 'local_g2_3')
// (7, 8, 'lutff_0/in_2')
// (7, 8, 'lutff_2/in_0')
// (7, 8, 'lutff_5/in_2')
// (7, 8, 'lutff_6/in_2')
// (7, 8, 'sp4_h_r_40')
// (7, 8, 'sp4_r_v_b_11')
// (8, 4, 'sp4_v_t_46')
// (8, 5, 'sp4_v_b_46')
// (8, 6, 'sp4_v_b_35')
// (8, 7, 'sp4_v_b_22')
// (8, 8, 'sp4_h_l_40')
// (8, 8, 'sp4_v_b_11')

wire n47;
// (0, 11, 'span12_horz_4')
// (1, 11, 'sp12_h_r_7')
// (2, 11, 'sp12_h_r_8')
// (3, 11, 'sp12_h_r_11')
// (4, 11, 'sp12_h_r_12')
// (5, 11, 'sp12_h_r_15')
// (6, 11, 'sp12_h_r_16')
// (7, 11, 'sp12_h_r_19')
// (7, 11, 'sp4_h_r_11')
// (8, 11, 'sp12_h_r_20')
// (8, 11, 'sp4_h_r_22')
// (9, 10, 'sp4_r_v_b_47')
// (9, 11, 'local_g0_7')
// (9, 11, 'local_g2_2')
// (9, 11, 'lutff_0/in_3')
// (9, 11, 'lutff_1/in_3')
// (9, 11, 'sp12_h_r_23')
// (9, 11, 'sp4_h_r_35')
// (9, 11, 'sp4_r_v_b_34')
// (9, 12, 'sp4_r_v_b_23')
// (9, 13, 'sp4_r_v_b_10')
// (10, 8, 'sp4_r_v_b_40')
// (10, 8, 'sp4_r_v_b_46')
// (10, 9, 'sp4_r_v_b_29')
// (10, 9, 'sp4_r_v_b_35')
// (10, 9, 'sp4_v_t_47')
// (10, 10, 'sp4_r_v_b_16')
// (10, 10, 'sp4_r_v_b_22')
// (10, 10, 'sp4_v_b_47')
// (10, 11, 'sp12_h_l_23')
// (10, 11, 'sp12_v_t_23')
// (10, 11, 'sp4_h_r_46')
// (10, 11, 'sp4_r_v_b_11')
// (10, 11, 'sp4_r_v_b_5')
// (10, 11, 'sp4_v_b_34')
// (10, 12, 'sp12_v_b_23')
// (10, 12, 'sp4_v_b_23')
// (10, 13, 'sp12_v_b_20')
// (10, 13, 'sp4_v_b_10')
// (10, 14, 'sp12_v_b_19')
// (10, 15, 'sp12_v_b_16')
// (10, 16, 'sp12_v_b_15')
// (10, 17, 'span12_vert_12')
// (11, 7, 'sp4_v_t_40')
// (11, 7, 'sp4_v_t_46')
// (11, 8, 'sp4_v_b_40')
// (11, 8, 'sp4_v_b_46')
// (11, 9, 'sp4_v_b_29')
// (11, 9, 'sp4_v_b_35')
// (11, 10, 'local_g0_6')
// (11, 10, 'local_g1_0')
// (11, 10, 'lutff_4/in_3')
// (11, 10, 'lutff_5/in_3')
// (11, 10, 'sp4_v_b_16')
// (11, 10, 'sp4_v_b_22')
// (11, 11, 'sp4_h_l_46')
// (11, 11, 'sp4_v_b_11')
// (11, 11, 'sp4_v_b_5')

wire n48;
// (0, 11, 'span12_horz_5')
// (1, 4, 'sp4_r_v_b_40')
// (1, 5, 'sp4_r_v_b_29')
// (1, 6, 'sp4_r_v_b_16')
// (1, 7, 'sp4_r_v_b_5')
// (1, 8, 'sp4_r_v_b_44')
// (1, 9, 'sp4_r_v_b_33')
// (1, 10, 'sp4_r_v_b_20')
// (1, 11, 'sp12_h_r_6')
// (1, 11, 'sp4_r_v_b_9')
// (2, 3, 'sp4_v_t_40')
// (2, 4, 'sp4_v_b_40')
// (2, 5, 'sp4_v_b_29')
// (2, 6, 'local_g0_0')
// (2, 6, 'lutff_6/in_0')
// (2, 6, 'sp4_v_b_16')
// (2, 7, 'sp4_v_b_5')
// (2, 7, 'sp4_v_t_44')
// (2, 8, 'sp4_v_b_44')
// (2, 9, 'sp4_v_b_33')
// (2, 10, 'sp4_v_b_20')
// (2, 11, 'sp12_h_r_9')
// (2, 11, 'sp4_h_r_4')
// (2, 11, 'sp4_v_b_9')
// (3, 11, 'sp12_h_r_10')
// (3, 11, 'sp4_h_r_17')
// (4, 11, 'sp12_h_r_13')
// (4, 11, 'sp4_h_r_28')
// (5, 11, 'sp12_h_r_14')
// (5, 11, 'sp4_h_r_41')
// (6, 10, 'neigh_op_tnr_5')
// (6, 11, 'neigh_op_rgt_5')
// (6, 11, 'sp12_h_r_17')
// (6, 11, 'sp4_h_l_41')
// (6, 12, 'neigh_op_bnr_5')
// (7, 10, 'local_g0_5')
// (7, 10, 'lutff_7/in_2')
// (7, 10, 'neigh_op_top_5')
// (7, 11, 'lutff_5/out')
// (7, 11, 'sp12_h_r_18')
// (7, 12, 'neigh_op_bot_5')
// (8, 10, 'neigh_op_tnl_5')
// (8, 11, 'local_g1_5')
// (8, 11, 'lutff_2/in_2')
// (8, 11, 'neigh_op_lft_5')
// (8, 11, 'sp12_h_r_21')
// (8, 12, 'neigh_op_bnl_5')
// (9, 11, 'sp12_h_r_22')
// (10, 11, 'sp12_h_l_22')

reg n49 = 0;
// (0, 11, 'span12_horz_8')
// (1, 10, 'neigh_op_tnr_2')
// (1, 11, 'neigh_op_rgt_2')
// (1, 11, 'sp12_h_r_11')
// (1, 12, 'neigh_op_bnr_2')
// (2, 10, 'neigh_op_top_2')
// (2, 11, 'lutff_2/out')
// (2, 11, 'sp12_h_r_12')
// (2, 12, 'neigh_op_bot_2')
// (3, 10, 'neigh_op_tnl_2')
// (3, 11, 'neigh_op_lft_2')
// (3, 11, 'sp12_h_r_15')
// (3, 12, 'neigh_op_bnl_2')
// (4, 11, 'sp12_h_r_16')
// (5, 11, 'local_g1_3')
// (5, 11, 'lutff_7/in_1')
// (5, 11, 'sp12_h_r_19')
// (6, 11, 'sp12_h_r_20')
// (7, 11, 'sp12_h_r_23')
// (8, 11, 'sp12_h_l_23')

reg n50 = 0;
// (0, 12, 'span12_horz_8')
// (1, 11, 'neigh_op_tnr_2')
// (1, 12, 'neigh_op_rgt_2')
// (1, 12, 'sp12_h_r_11')
// (1, 13, 'neigh_op_bnr_2')
// (2, 11, 'neigh_op_top_2')
// (2, 12, 'lutff_2/out')
// (2, 12, 'sp12_h_r_12')
// (2, 13, 'neigh_op_bot_2')
// (3, 11, 'neigh_op_tnl_2')
// (3, 12, 'neigh_op_lft_2')
// (3, 12, 'sp12_h_r_15')
// (3, 13, 'neigh_op_bnl_2')
// (4, 12, 'local_g0_0')
// (4, 12, 'lutff_2/in_0')
// (4, 12, 'sp12_h_r_16')
// (5, 12, 'sp12_h_r_19')
// (6, 12, 'sp12_h_r_20')
// (7, 12, 'sp12_h_r_23')
// (8, 12, 'sp12_h_l_23')

reg n51 = 0;
// (0, 13, 'span12_horz_12')
// (1, 12, 'neigh_op_tnr_4')
// (1, 13, 'neigh_op_rgt_4')
// (1, 13, 'sp12_h_r_15')
// (1, 13, 'sp4_h_r_9')
// (1, 14, 'neigh_op_bnr_4')
// (2, 12, 'neigh_op_top_4')
// (2, 13, 'lutff_4/out')
// (2, 13, 'sp12_h_r_16')
// (2, 13, 'sp4_h_r_20')
// (2, 14, 'neigh_op_bot_4')
// (3, 12, 'neigh_op_tnl_4')
// (3, 13, 'neigh_op_lft_4')
// (3, 13, 'sp12_h_r_19')
// (3, 13, 'sp4_h_r_33')
// (3, 14, 'neigh_op_bnl_4')
// (4, 10, 'sp4_r_v_b_38')
// (4, 11, 'sp4_r_v_b_27')
// (4, 12, 'sp4_r_v_b_14')
// (4, 13, 'local_g1_4')
// (4, 13, 'lutff_5/in_0')
// (4, 13, 'sp12_h_r_20')
// (4, 13, 'sp4_h_r_44')
// (4, 13, 'sp4_r_v_b_3')
// (5, 9, 'sp4_v_t_38')
// (5, 10, 'sp4_v_b_38')
// (5, 11, 'sp4_v_b_27')
// (5, 12, 'local_g1_6')
// (5, 12, 'lutff_3/in_0')
// (5, 12, 'lutff_5/in_0')
// (5, 12, 'sp4_v_b_14')
// (5, 13, 'local_g1_7')
// (5, 13, 'lutff_2/in_0')
// (5, 13, 'sp12_h_r_23')
// (5, 13, 'sp4_h_l_44')
// (5, 13, 'sp4_v_b_3')
// (6, 13, 'sp12_h_l_23')

wire rst;
// (0, 14, 'io_1/D_IN_0')
// (0, 14, 'io_1/PAD')
// (0, 14, 'span4_horz_28')
// (1, 3, 'sp4_r_v_b_37')
// (1, 4, 'sp4_r_v_b_24')
// (1, 5, 'sp4_r_v_b_13')
// (1, 6, 'sp4_r_v_b_0')
// (1, 7, 'sp4_r_v_b_37')
// (1, 8, 'sp4_r_v_b_24')
// (1, 9, 'sp4_r_v_b_13')
// (1, 10, 'sp4_r_v_b_0')
// (1, 11, 'sp4_r_v_b_41')
// (1, 12, 'local_g0_4')
// (1, 12, 'lutff_5/in_3')
// (1, 12, 'sp4_r_v_b_28')
// (1, 13, 'neigh_op_tnl_2')
// (1, 13, 'neigh_op_tnl_6')
// (1, 13, 'sp4_r_v_b_17')
// (1, 14, 'neigh_op_lft_2')
// (1, 14, 'neigh_op_lft_6')
// (1, 14, 'sp4_h_r_41')
// (1, 14, 'sp4_r_v_b_4')
// (1, 15, 'neigh_op_bnl_2')
// (1, 15, 'neigh_op_bnl_6')
// (2, 2, 'sp4_v_t_37')
// (2, 3, 'sp4_v_b_37')
// (2, 4, 'local_g2_0')
// (2, 4, 'lutff_1/in_3')
// (2, 4, 'sp4_v_b_24')
// (2, 5, 'sp4_v_b_13')
// (2, 6, 'sp4_h_r_5')
// (2, 6, 'sp4_v_b_0')
// (2, 6, 'sp4_v_t_37')
// (2, 7, 'sp4_v_b_37')
// (2, 8, 'sp4_v_b_24')
// (2, 9, 'sp4_v_b_13')
// (2, 10, 'sp4_v_b_0')
// (2, 10, 'sp4_v_t_41')
// (2, 11, 'sp4_v_b_41')
// (2, 12, 'sp4_v_b_28')
// (2, 13, 'sp4_v_b_17')
// (2, 14, 'sp4_h_l_41')
// (2, 14, 'sp4_v_b_4')
// (3, 6, 'sp4_h_r_16')
// (4, 6, 'sp4_h_r_29')
// (5, 6, 'sp4_h_r_40')
// (6, 6, 'sp4_h_l_40')
// (6, 6, 'sp4_h_r_1')
// (6, 6, 'sp4_h_r_5')
// (7, 3, 'local_g3_2')
// (7, 3, 'lutff_2/in_3')
// (7, 3, 'sp4_r_v_b_42')
// (7, 4, 'sp4_r_v_b_31')
// (7, 5, 'sp4_r_v_b_18')
// (7, 6, 'sp4_h_r_12')
// (7, 6, 'sp4_h_r_16')
// (7, 6, 'sp4_r_v_b_7')
// (8, 2, 'sp4_h_r_1')
// (8, 2, 'sp4_v_t_42')
// (8, 3, 'sp4_v_b_42')
// (8, 4, 'sp4_v_b_31')
// (8, 5, 'sp4_v_b_18')
// (8, 6, 'sp4_h_r_25')
// (8, 6, 'sp4_h_r_29')
// (8, 6, 'sp4_v_b_7')
// (9, 2, 'sp4_h_r_12')
// (9, 3, 'local_g2_4')
// (9, 3, 'lutff_5/in_1')
// (9, 3, 'sp4_r_v_b_36')
// (9, 3, 'sp4_r_v_b_40')
// (9, 4, 'local_g0_5')
// (9, 4, 'local_g1_5')
// (9, 4, 'lutff_4/in_3')
// (9, 4, 'lutff_5/in_3')
// (9, 4, 'lutff_7/in_1')
// (9, 4, 'sp4_r_v_b_25')
// (9, 4, 'sp4_r_v_b_29')
// (9, 5, 'sp4_r_v_b_12')
// (9, 5, 'sp4_r_v_b_16')
// (9, 6, 'local_g2_0')
// (9, 6, 'lutff_1/in_3')
// (9, 6, 'sp4_h_r_36')
// (9, 6, 'sp4_h_r_40')
// (9, 6, 'sp4_r_v_b_1')
// (9, 6, 'sp4_r_v_b_5')
// (10, 2, 'sp4_h_r_1')
// (10, 2, 'sp4_h_r_25')
// (10, 2, 'sp4_v_t_36')
// (10, 2, 'sp4_v_t_40')
// (10, 3, 'sp4_v_b_36')
// (10, 3, 'sp4_v_b_40')
// (10, 4, 'sp4_v_b_25')
// (10, 4, 'sp4_v_b_29')
// (10, 5, 'sp4_v_b_12')
// (10, 5, 'sp4_v_b_16')
// (10, 6, 'sp4_h_l_36')
// (10, 6, 'sp4_h_l_40')
// (10, 6, 'sp4_v_b_1')
// (10, 6, 'sp4_v_b_5')
// (11, 2, 'sp4_h_r_12')
// (11, 2, 'sp4_h_r_36')
// (11, 3, 'local_g2_4')
// (11, 3, 'lutff_global/s_r')
// (11, 3, 'sp4_r_v_b_36')
// (11, 4, 'local_g1_1')
// (11, 4, 'lutff_7/in_3')
// (11, 4, 'sp4_r_v_b_25')
// (11, 5, 'local_g2_4')
// (11, 5, 'lutff_1/in_3')
// (11, 5, 'sp4_r_v_b_12')
// (11, 6, 'sp4_r_v_b_1')
// (12, 2, 'sp4_h_l_36')
// (12, 2, 'sp4_h_r_1')
// (12, 2, 'sp4_h_r_25')
// (12, 2, 'sp4_v_t_36')
// (12, 3, 'sp4_v_b_36')
// (12, 4, 'sp4_v_b_25')
// (12, 5, 'sp4_v_b_12')
// (12, 6, 'sp4_v_b_1')
// (13, 2, 'span4_horz_1')
// (13, 2, 'span4_horz_25')

reg n53 = 0;
// (0, 14, 'span12_horz_12')
// (1, 13, 'neigh_op_tnr_4')
// (1, 14, 'neigh_op_rgt_4')
// (1, 14, 'sp12_h_r_15')
// (1, 15, 'neigh_op_bnr_4')
// (2, 13, 'neigh_op_top_4')
// (2, 14, 'lutff_4/out')
// (2, 14, 'sp12_h_r_16')
// (2, 15, 'neigh_op_bot_4')
// (3, 13, 'neigh_op_tnl_4')
// (3, 14, 'neigh_op_lft_4')
// (3, 14, 'sp12_h_r_19')
// (3, 15, 'neigh_op_bnl_4')
// (4, 14, 'local_g0_4')
// (4, 14, 'lutff_6/in_0')
// (4, 14, 'sp12_h_r_20')
// (5, 9, 'sp4_r_v_b_39')
// (5, 10, 'local_g1_2')
// (5, 10, 'lutff_3/in_0')
// (5, 10, 'sp4_r_v_b_26')
// (5, 11, 'sp4_r_v_b_15')
// (5, 12, 'local_g1_2')
// (5, 12, 'lutff_1/in_0')
// (5, 12, 'sp4_r_v_b_2')
// (5, 14, 'local_g0_7')
// (5, 14, 'lutff_5/in_0')
// (5, 14, 'sp12_h_r_23')
// (6, 2, 'sp12_v_t_23')
// (6, 3, 'sp12_v_b_23')
// (6, 4, 'sp12_v_b_20')
// (6, 5, 'sp12_v_b_19')
// (6, 6, 'sp12_v_b_16')
// (6, 7, 'sp12_v_b_15')
// (6, 8, 'sp12_v_b_12')
// (6, 8, 'sp4_v_t_39')
// (6, 9, 'sp12_v_b_11')
// (6, 9, 'sp4_v_b_39')
// (6, 10, 'sp12_v_b_8')
// (6, 10, 'sp4_v_b_26')
// (6, 11, 'sp12_v_b_7')
// (6, 11, 'sp4_v_b_15')
// (6, 12, 'sp12_v_b_4')
// (6, 12, 'sp4_v_b_2')
// (6, 13, 'sp12_v_b_3')
// (6, 14, 'sp12_h_l_23')
// (6, 14, 'sp12_v_b_0')

reg n54 = 0;
// (0, 14, 'span12_horz_2')
// (1, 14, 'sp12_h_r_5')
// (2, 14, 'local_g0_6')
// (2, 14, 'lutff_2/in_0')
// (2, 14, 'sp12_h_r_6')
// (3, 13, 'neigh_op_tnr_1')
// (3, 14, 'neigh_op_rgt_1')
// (3, 14, 'sp12_h_r_9')
// (3, 15, 'neigh_op_bnr_1')
// (4, 13, 'neigh_op_top_1')
// (4, 14, 'lutff_1/out')
// (4, 14, 'sp12_h_r_10')
// (4, 15, 'neigh_op_bot_1')
// (5, 13, 'neigh_op_tnl_1')
// (5, 14, 'neigh_op_lft_1')
// (5, 14, 'sp12_h_r_13')
// (5, 15, 'neigh_op_bnl_1')
// (6, 14, 'sp12_h_r_14')
// (7, 14, 'sp12_h_r_17')
// (8, 14, 'sp12_h_r_18')
// (9, 14, 'sp12_h_r_21')
// (10, 14, 'sp12_h_r_22')
// (11, 14, 'sp12_h_l_22')

wire n55;
// (1, 1, 'neigh_op_tnr_0')
// (1, 1, 'sp4_r_v_b_45')
// (1, 2, 'neigh_op_rgt_0')
// (1, 2, 'sp4_r_v_b_32')
// (1, 3, 'neigh_op_bnr_0')
// (1, 3, 'sp4_r_v_b_21')
// (1, 4, 'sp4_r_v_b_8')
// (2, 0, 'span4_vert_45')
// (2, 1, 'neigh_op_top_0')
// (2, 1, 'sp4_v_b_45')
// (2, 2, 'lutff_0/out')
// (2, 2, 'sp4_v_b_32')
// (2, 3, 'neigh_op_bot_0')
// (2, 3, 'sp4_v_b_21')
// (2, 4, 'local_g1_0')
// (2, 4, 'lutff_1/in_2')
// (2, 4, 'sp4_v_b_8')
// (3, 1, 'neigh_op_tnl_0')
// (3, 2, 'neigh_op_lft_0')
// (3, 3, 'neigh_op_bnl_0')

wire n56;
// (1, 1, 'neigh_op_tnr_4')
// (1, 2, 'neigh_op_rgt_4')
// (1, 3, 'neigh_op_bnr_4')
// (2, 1, 'neigh_op_top_4')
// (2, 2, 'lutff_4/out')
// (2, 2, 'sp4_h_r_8')
// (2, 3, 'neigh_op_bot_4')
// (3, 1, 'neigh_op_tnl_4')
// (3, 2, 'neigh_op_lft_4')
// (3, 2, 'sp4_h_r_21')
// (3, 3, 'neigh_op_bnl_4')
// (4, 2, 'sp4_h_r_32')
// (5, 2, 'sp4_h_r_45')
// (5, 3, 'local_g2_4')
// (5, 3, 'lutff_2/in_2')
// (5, 3, 'sp4_r_v_b_36')
// (5, 4, 'sp4_r_v_b_25')
// (5, 5, 'sp4_r_v_b_12')
// (5, 6, 'sp4_r_v_b_1')
// (6, 2, 'sp4_h_l_45')
// (6, 2, 'sp4_v_t_36')
// (6, 3, 'sp4_v_b_36')
// (6, 4, 'sp4_v_b_25')
// (6, 5, 'sp4_v_b_12')
// (6, 6, 'sp4_v_b_1')

reg n57 = 0;
// (1, 2, 'neigh_op_tnr_2')
// (1, 3, 'neigh_op_rgt_2')
// (1, 3, 'sp4_r_v_b_36')
// (1, 4, 'neigh_op_bnr_2')
// (1, 4, 'sp4_r_v_b_25')
// (1, 5, 'sp4_r_v_b_12')
// (1, 6, 'sp4_r_v_b_1')
// (2, 2, 'neigh_op_top_2')
// (2, 2, 'sp4_v_t_36')
// (2, 3, 'local_g0_2')
// (2, 3, 'lutff_2/in_2')
// (2, 3, 'lutff_2/out')
// (2, 3, 'sp4_v_b_36')
// (2, 4, 'local_g1_2')
// (2, 4, 'lutff_3/in_2')
// (2, 4, 'neigh_op_bot_2')
// (2, 4, 'sp4_v_b_25')
// (2, 5, 'local_g1_4')
// (2, 5, 'lutff_3/in_2')
// (2, 5, 'sp4_v_b_12')
// (2, 6, 'sp4_v_b_1')
// (3, 2, 'neigh_op_tnl_2')
// (3, 3, 'neigh_op_lft_2')
// (3, 4, 'neigh_op_bnl_2')

reg n58 = 0;
// (1, 2, 'neigh_op_tnr_3')
// (1, 3, 'neigh_op_rgt_3')
// (1, 4, 'neigh_op_bnr_3')
// (2, 2, 'neigh_op_top_3')
// (2, 3, 'local_g0_3')
// (2, 3, 'lutff_3/in_2')
// (2, 3, 'lutff_3/out')
// (2, 3, 'sp4_r_v_b_39')
// (2, 4, 'local_g0_2')
// (2, 4, 'lutff_3/in_1')
// (2, 4, 'neigh_op_bot_3')
// (2, 4, 'sp4_r_v_b_26')
// (2, 5, 'local_g2_7')
// (2, 5, 'lutff_2/in_1')
// (2, 5, 'lutff_3/in_0')
// (2, 5, 'sp4_r_v_b_15')
// (2, 6, 'sp4_r_v_b_2')
// (3, 2, 'neigh_op_tnl_3')
// (3, 2, 'sp4_v_t_39')
// (3, 3, 'neigh_op_lft_3')
// (3, 3, 'sp4_v_b_39')
// (3, 4, 'neigh_op_bnl_3')
// (3, 4, 'sp4_v_b_26')
// (3, 5, 'sp4_v_b_15')
// (3, 6, 'sp4_v_b_2')

reg n59 = 0;
// (1, 2, 'neigh_op_tnr_6')
// (1, 3, 'neigh_op_rgt_6')
// (1, 3, 'sp4_h_r_1')
// (1, 4, 'neigh_op_bnr_6')
// (2, 2, 'local_g0_6')
// (2, 2, 'lutff_4/in_0')
// (2, 2, 'neigh_op_top_6')
// (2, 3, 'local_g0_6')
// (2, 3, 'lutff_6/in_2')
// (2, 3, 'lutff_6/out')
// (2, 3, 'sp4_h_r_12')
// (2, 4, 'neigh_op_bot_6')
// (3, 2, 'neigh_op_tnl_6')
// (3, 3, 'neigh_op_lft_6')
// (3, 3, 'sp4_h_r_25')
// (3, 4, 'neigh_op_bnl_6')
// (4, 1, 'sp4_r_v_b_24')
// (4, 1, 'sp4_r_v_b_25')
// (4, 1, 'sp4_r_v_b_29')
// (4, 1, 'sp4_r_v_b_31')
// (4, 2, 'sp4_r_v_b_12')
// (4, 2, 'sp4_r_v_b_13')
// (4, 2, 'sp4_r_v_b_16')
// (4, 2, 'sp4_r_v_b_18')
// (4, 3, 'local_g2_4')
// (4, 3, 'lutff_5/in_3')
// (4, 3, 'sp4_h_r_36')
// (4, 3, 'sp4_r_v_b_0')
// (4, 3, 'sp4_r_v_b_1')
// (4, 3, 'sp4_r_v_b_5')
// (4, 3, 'sp4_r_v_b_7')
// (4, 4, 'sp4_r_v_b_44')
// (4, 5, 'sp4_r_v_b_33')
// (4, 6, 'sp4_r_v_b_20')
// (4, 7, 'sp4_r_v_b_9')
// (5, 0, 'span4_vert_24')
// (5, 0, 'span4_vert_25')
// (5, 0, 'span4_vert_29')
// (5, 0, 'span4_vert_31')
// (5, 1, 'sp4_v_b_24')
// (5, 1, 'sp4_v_b_25')
// (5, 1, 'sp4_v_b_29')
// (5, 1, 'sp4_v_b_31')
// (5, 2, 'local_g0_0')
// (5, 2, 'local_g1_2')
// (5, 2, 'lutff_3/in_2')
// (5, 2, 'lutff_4/in_2')
// (5, 2, 'sp4_v_b_12')
// (5, 2, 'sp4_v_b_13')
// (5, 2, 'sp4_v_b_16')
// (5, 2, 'sp4_v_b_18')
// (5, 3, 'local_g0_0')
// (5, 3, 'local_g0_1')
// (5, 3, 'lutff_0/in_0')
// (5, 3, 'lutff_1/in_0')
// (5, 3, 'lutff_3/in_2')
// (5, 3, 'sp4_h_l_36')
// (5, 3, 'sp4_v_b_0')
// (5, 3, 'sp4_v_b_1')
// (5, 3, 'sp4_v_b_5')
// (5, 3, 'sp4_v_b_7')
// (5, 3, 'sp4_v_t_44')
// (5, 4, 'sp4_v_b_44')
// (5, 5, 'sp4_v_b_33')
// (5, 6, 'sp4_v_b_20')
// (5, 7, 'sp4_v_b_9')

wire n60;
// (1, 3, 'neigh_op_tnr_1')
// (1, 4, 'neigh_op_rgt_1')
// (1, 5, 'neigh_op_bnr_1')
// (1, 9, 'sp4_r_v_b_38')
// (1, 10, 'sp4_r_v_b_27')
// (1, 11, 'sp4_r_v_b_14')
// (1, 12, 'local_g1_3')
// (1, 12, 'lutff_global/cen')
// (1, 12, 'sp4_r_v_b_3')
// (2, 1, 'sp12_v_t_22')
// (2, 2, 'sp12_v_b_22')
// (2, 3, 'neigh_op_top_1')
// (2, 3, 'sp12_v_b_21')
// (2, 4, 'lutff_1/out')
// (2, 4, 'sp12_v_b_18')
// (2, 5, 'neigh_op_bot_1')
// (2, 5, 'sp12_v_b_17')
// (2, 6, 'sp12_v_b_14')
// (2, 7, 'sp12_v_b_13')
// (2, 8, 'sp12_v_b_10')
// (2, 8, 'sp4_v_t_38')
// (2, 9, 'sp12_v_b_9')
// (2, 9, 'sp4_v_b_38')
// (2, 10, 'sp12_v_b_6')
// (2, 10, 'sp4_v_b_27')
// (2, 11, 'sp12_v_b_5')
// (2, 11, 'sp4_v_b_14')
// (2, 12, 'sp12_v_b_2')
// (2, 12, 'sp4_v_b_3')
// (2, 13, 'sp12_v_b_1')
// (3, 3, 'neigh_op_tnl_1')
// (3, 4, 'neigh_op_lft_1')
// (3, 5, 'neigh_op_bnl_1')

wire n61;
// (1, 3, 'neigh_op_tnr_3')
// (1, 4, 'neigh_op_rgt_3')
// (1, 5, 'neigh_op_bnr_3')
// (2, 3, 'neigh_op_top_3')
// (2, 4, 'local_g1_3')
// (2, 4, 'lutff_1/in_1')
// (2, 4, 'lutff_3/out')
// (2, 5, 'neigh_op_bot_3')
// (3, 3, 'neigh_op_tnl_3')
// (3, 4, 'neigh_op_lft_3')
// (3, 5, 'neigh_op_bnl_3')

reg n62 = 0;
// (1, 3, 'neigh_op_tnr_6')
// (1, 4, 'neigh_op_rgt_6')
// (1, 5, 'neigh_op_bnr_6')
// (2, 3, 'local_g1_6')
// (2, 3, 'lutff_0/in_1')
// (2, 3, 'neigh_op_top_6')
// (2, 4, 'local_g0_6')
// (2, 4, 'local_g1_6')
// (2, 4, 'lutff_3/in_3')
// (2, 4, 'lutff_6/in_3')
// (2, 4, 'lutff_6/out')
// (2, 4, 'lutff_7/in_3')
// (2, 5, 'local_g0_6')
// (2, 5, 'local_g1_6')
// (2, 5, 'lutff_0/in_3')
// (2, 5, 'lutff_2/in_3')
// (2, 5, 'lutff_3/in_3')
// (2, 5, 'neigh_op_bot_6')
// (3, 3, 'neigh_op_tnl_6')
// (3, 4, 'neigh_op_lft_6')
// (3, 5, 'neigh_op_bnl_6')

reg n63 = 0;
// (1, 3, 'neigh_op_tnr_7')
// (1, 4, 'neigh_op_rgt_7')
// (1, 5, 'neigh_op_bnr_7')
// (2, 3, 'local_g0_7')
// (2, 3, 'lutff_1/in_2')
// (2, 3, 'neigh_op_top_7')
// (2, 4, 'local_g0_7')
// (2, 4, 'lutff_3/in_0')
// (2, 4, 'lutff_7/in_2')
// (2, 4, 'lutff_7/out')
// (2, 5, 'local_g1_7')
// (2, 5, 'lutff_0/in_2')
// (2, 5, 'lutff_2/in_2')
// (2, 5, 'lutff_3/in_1')
// (2, 5, 'neigh_op_bot_7')
// (3, 3, 'neigh_op_tnl_7')
// (3, 4, 'neigh_op_lft_7')
// (3, 5, 'neigh_op_bnl_7')

wire n64;
// (1, 3, 'sp12_h_r_0')
// (2, 3, 'sp12_h_r_3')
// (3, 3, 'sp12_h_r_4')
// (4, 2, 'neigh_op_tnr_0')
// (4, 3, 'neigh_op_rgt_0')
// (4, 3, 'sp12_h_r_7')
// (4, 4, 'neigh_op_bnr_0')
// (5, 2, 'neigh_op_top_0')
// (5, 3, 'lutff_0/out')
// (5, 3, 'sp12_h_r_8')
// (5, 4, 'neigh_op_bot_0')
// (6, 2, 'neigh_op_tnl_0')
// (6, 3, 'neigh_op_lft_0')
// (6, 3, 'sp12_h_r_11')
// (6, 4, 'neigh_op_bnl_0')
// (7, 3, 'local_g0_4')
// (7, 3, 'lutff_2/in_2')
// (7, 3, 'sp12_h_r_12')
// (8, 3, 'sp12_h_r_15')
// (9, 3, 'sp12_h_r_16')
// (10, 3, 'sp12_h_r_19')
// (11, 3, 'sp12_h_r_20')
// (12, 3, 'sp12_h_r_23')
// (13, 3, 'span12_horz_23')

wire n65;
// (1, 4, 'neigh_op_tnr_0')
// (1, 5, 'neigh_op_rgt_0')
// (1, 6, 'neigh_op_bnr_0')
// (2, 3, 'sp4_r_v_b_41')
// (2, 4, 'neigh_op_top_0')
// (2, 4, 'sp4_r_v_b_28')
// (2, 5, 'local_g1_0')
// (2, 5, 'lutff_0/out')
// (2, 5, 'lutff_1/in_0')
// (2, 5, 'sp4_r_v_b_17')
// (2, 6, 'neigh_op_bot_0')
// (2, 6, 'sp4_r_v_b_4')
// (3, 2, 'sp4_v_t_41')
// (3, 3, 'sp4_v_b_41')
// (3, 4, 'neigh_op_tnl_0')
// (3, 4, 'sp4_v_b_28')
// (3, 5, 'neigh_op_lft_0')
// (3, 5, 'sp4_v_b_17')
// (3, 6, 'neigh_op_bnl_0')
// (3, 6, 'sp4_h_r_10')
// (3, 6, 'sp4_v_b_4')
// (4, 6, 'local_g1_7')
// (4, 6, 'lutff_5/in_3')
// (4, 6, 'sp4_h_r_23')
// (5, 6, 'sp4_h_r_34')
// (6, 6, 'sp4_h_r_47')
// (7, 6, 'sp4_h_l_47')

reg n66 = 0;
// (1, 5, 'sp4_h_r_1')
// (2, 5, 'local_g0_4')
// (2, 5, 'lutff_global/s_r')
// (2, 5, 'sp4_h_r_12')
// (3, 5, 'sp4_h_r_25')
// (4, 5, 'sp4_h_r_36')
// (5, 5, 'sp4_h_l_36')
// (5, 5, 'sp4_h_r_1')
// (6, 5, 'sp4_h_r_12')
// (7, 5, 'sp4_h_r_25')
// (8, 2, 'sp4_r_v_b_38')
// (8, 3, 'sp4_r_v_b_27')
// (8, 4, 'sp4_r_v_b_14')
// (8, 5, 'sp4_h_r_36')
// (8, 5, 'sp4_r_v_b_3')
// (9, 1, 'sp4_v_t_38')
// (9, 2, 'sp4_v_b_38')
// (9, 3, 'local_g2_3')
// (9, 3, 'lutff_5/in_2')
// (9, 3, 'sp4_v_b_27')
// (9, 4, 'sp4_v_b_14')
// (9, 5, 'local_g0_2')
// (9, 5, 'lutff_1/in_1')
// (9, 5, 'sp4_h_l_36')
// (9, 5, 'sp4_h_r_10')
// (9, 5, 'sp4_v_b_3')
// (10, 4, 'neigh_op_tnr_1')
// (10, 5, 'neigh_op_rgt_1')
// (10, 5, 'sp4_h_r_23')
// (10, 6, 'neigh_op_bnr_1')
// (11, 2, 'sp4_r_v_b_38')
// (11, 3, 'local_g1_3')
// (11, 3, 'lutff_7/in_1')
// (11, 3, 'sp4_r_v_b_27')
// (11, 4, 'local_g0_1')
// (11, 4, 'lutff_1/in_0')
// (11, 4, 'neigh_op_top_1')
// (11, 4, 'sp4_r_v_b_14')
// (11, 5, 'local_g0_1')
// (11, 5, 'lutff_1/in_2')
// (11, 5, 'lutff_1/out')
// (11, 5, 'sp4_h_r_34')
// (11, 5, 'sp4_r_v_b_3')
// (11, 6, 'neigh_op_bot_1')
// (12, 1, 'sp4_v_t_38')
// (12, 2, 'sp4_v_b_38')
// (12, 3, 'sp4_v_b_27')
// (12, 4, 'neigh_op_tnl_1')
// (12, 4, 'sp4_v_b_14')
// (12, 5, 'neigh_op_lft_1')
// (12, 5, 'sp4_h_r_47')
// (12, 5, 'sp4_v_b_3')
// (12, 6, 'neigh_op_bnl_1')
// (13, 5, 'span4_horz_47')

wire n67;
// (1, 5, 'sp4_h_r_5')
// (2, 5, 'sp4_h_r_16')
// (3, 5, 'sp4_h_r_29')
// (4, 2, 'neigh_op_tnr_4')
// (4, 2, 'sp4_r_v_b_37')
// (4, 3, 'neigh_op_rgt_4')
// (4, 3, 'sp4_r_v_b_24')
// (4, 4, 'neigh_op_bnr_4')
// (4, 4, 'sp4_r_v_b_13')
// (4, 5, 'local_g1_0')
// (4, 5, 'local_g2_0')
// (4, 5, 'lutff_3/in_1')
// (4, 5, 'lutff_4/in_1')
// (4, 5, 'sp4_h_r_40')
// (4, 5, 'sp4_r_v_b_0')
// (5, 1, 'sp4_v_t_37')
// (5, 2, 'neigh_op_top_4')
// (5, 2, 'sp4_v_b_37')
// (5, 3, 'lutff_4/out')
// (5, 3, 'sp4_v_b_24')
// (5, 4, 'neigh_op_bot_4')
// (5, 4, 'sp4_v_b_13')
// (5, 5, 'local_g1_0')
// (5, 5, 'lutff_7/in_2')
// (5, 5, 'sp4_h_l_40')
// (5, 5, 'sp4_v_b_0')
// (6, 2, 'neigh_op_tnl_4')
// (6, 3, 'neigh_op_lft_4')
// (6, 4, 'neigh_op_bnl_4')

wire n68;
// (1, 6, 'sp12_h_r_0')
// (2, 6, 'sp12_h_r_3')
// (3, 6, 'sp12_h_r_4')
// (4, 6, 'sp12_h_r_7')
// (5, 6, 'local_g0_0')
// (5, 6, 'local_g1_0')
// (5, 6, 'lutff_1/in_1')
// (5, 6, 'lutff_4/in_3')
// (5, 6, 'sp12_h_r_8')
// (6, 5, 'neigh_op_tnr_2')
// (6, 6, 'local_g2_2')
// (6, 6, 'local_g3_2')
// (6, 6, 'lutff_0/in_2')
// (6, 6, 'lutff_3/in_1')
// (6, 6, 'lutff_6/in_1')
// (6, 6, 'neigh_op_rgt_2')
// (6, 6, 'sp12_h_r_11')
// (6, 7, 'neigh_op_bnr_2')
// (7, 5, 'neigh_op_top_2')
// (7, 6, 'local_g1_2')
// (7, 6, 'lutff_1/in_0')
// (7, 6, 'lutff_2/out')
// (7, 6, 'lutff_6/in_3')
// (7, 6, 'sp12_h_r_12')
// (7, 7, 'neigh_op_bot_2')
// (8, 5, 'neigh_op_tnl_2')
// (8, 6, 'neigh_op_lft_2')
// (8, 6, 'sp12_h_r_15')
// (8, 7, 'neigh_op_bnl_2')
// (9, 6, 'sp12_h_r_16')
// (10, 6, 'sp12_h_r_19')
// (11, 6, 'sp12_h_r_20')
// (12, 6, 'sp12_h_r_23')
// (13, 6, 'span12_horz_23')

reg n69 = 0;
// (1, 6, 'sp12_h_r_1')
// (2, 6, 'sp12_h_r_2')
// (3, 5, 'neigh_op_tnr_7')
// (3, 6, 'neigh_op_rgt_7')
// (3, 6, 'sp12_h_r_5')
// (3, 7, 'neigh_op_bnr_7')
// (4, 5, 'neigh_op_top_7')
// (4, 6, 'local_g0_7')
// (4, 6, 'lutff_1/in_0')
// (4, 6, 'lutff_7/out')
// (4, 6, 'sp12_h_r_6')
// (4, 7, 'neigh_op_bot_7')
// (5, 5, 'neigh_op_tnl_7')
// (5, 6, 'neigh_op_lft_7')
// (5, 6, 'sp12_h_r_9')
// (5, 7, 'neigh_op_bnl_7')
// (6, 6, 'sp12_h_r_10')
// (7, 6, 'sp12_h_r_13')
// (8, 6, 'local_g1_6')
// (8, 6, 'lutff_4/in_3')
// (8, 6, 'sp12_h_r_14')
// (9, 6, 'sp12_h_r_17')
// (10, 6, 'sp12_h_r_18')
// (11, 6, 'sp12_h_r_21')
// (12, 6, 'sp12_h_r_22')
// (13, 6, 'span12_horz_22')

reg n70 = 0;
// (1, 6, 'sp4_r_v_b_41')
// (1, 7, 'sp4_r_v_b_28')
// (1, 8, 'neigh_op_tnr_2')
// (1, 8, 'sp4_r_v_b_17')
// (1, 9, 'neigh_op_rgt_2')
// (1, 9, 'sp4_r_v_b_4')
// (1, 10, 'neigh_op_bnr_2')
// (2, 5, 'sp4_v_t_41')
// (2, 6, 'sp4_v_b_41')
// (2, 7, 'sp4_v_b_28')
// (2, 8, 'local_g1_1')
// (2, 8, 'lutff_3/in_1')
// (2, 8, 'neigh_op_top_2')
// (2, 8, 'sp4_v_b_17')
// (2, 9, 'lutff_2/out')
// (2, 9, 'sp4_v_b_4')
// (2, 10, 'neigh_op_bot_2')
// (3, 8, 'neigh_op_tnl_2')
// (3, 9, 'neigh_op_lft_2')
// (3, 10, 'neigh_op_bnl_2')

reg n71 = 0;
// (1, 7, 'neigh_op_tnr_3')
// (1, 8, 'neigh_op_rgt_3')
// (1, 9, 'neigh_op_bnr_3')
// (2, 6, 'sp4_r_v_b_47')
// (2, 7, 'neigh_op_top_3')
// (2, 7, 'sp4_r_v_b_34')
// (2, 8, 'lutff_3/out')
// (2, 8, 'sp4_r_v_b_23')
// (2, 9, 'neigh_op_bot_3')
// (2, 9, 'sp4_r_v_b_10')
// (3, 5, 'sp4_v_t_47')
// (3, 6, 'sp4_v_b_47')
// (3, 7, 'neigh_op_tnl_3')
// (3, 7, 'sp4_v_b_34')
// (3, 8, 'neigh_op_lft_3')
// (3, 8, 'sp4_v_b_23')
// (3, 9, 'neigh_op_bnl_3')
// (3, 9, 'sp4_h_r_4')
// (3, 9, 'sp4_v_b_10')
// (4, 9, 'local_g0_1')
// (4, 9, 'lutff_6/in_1')
// (4, 9, 'sp4_h_r_17')
// (5, 9, 'sp4_h_r_28')
// (6, 9, 'sp4_h_r_41')
// (7, 9, 'sp4_h_l_41')

reg n72 = 0;
// (1, 7, 'neigh_op_tnr_7')
// (1, 8, 'neigh_op_rgt_7')
// (1, 9, 'neigh_op_bnr_7')
// (2, 7, 'neigh_op_top_7')
// (2, 8, 'local_g0_7')
// (2, 8, 'lutff_0/in_1')
// (2, 8, 'lutff_7/out')
// (2, 9, 'neigh_op_bot_7')
// (3, 7, 'neigh_op_tnl_7')
// (3, 8, 'neigh_op_lft_7')
// (3, 9, 'neigh_op_bnl_7')

reg n73 = 0;
// (1, 8, 'neigh_op_tnr_5')
// (1, 9, 'neigh_op_rgt_5')
// (1, 9, 'sp12_h_r_1')
// (1, 10, 'neigh_op_bnr_5')
// (2, 8, 'neigh_op_top_5')
// (2, 9, 'lutff_5/out')
// (2, 9, 'sp12_h_r_2')
// (2, 10, 'neigh_op_bot_5')
// (3, 8, 'neigh_op_tnl_5')
// (3, 9, 'neigh_op_lft_5')
// (3, 9, 'sp12_h_r_5')
// (3, 10, 'neigh_op_bnl_5')
// (4, 9, 'local_g1_6')
// (4, 9, 'lutff_0/in_1')
// (4, 9, 'sp12_h_r_6')
// (5, 9, 'sp12_h_r_9')
// (6, 9, 'sp12_h_r_10')
// (7, 9, 'sp12_h_r_13')
// (8, 9, 'sp12_h_r_14')
// (9, 9, 'sp12_h_r_17')
// (10, 9, 'sp12_h_r_18')
// (11, 9, 'sp12_h_r_21')
// (12, 9, 'sp12_h_r_22')
// (13, 9, 'span12_horz_22')

reg n74 = 0;
// (1, 8, 'sp4_h_r_7')
// (2, 8, 'local_g0_2')
// (2, 8, 'lutff_0/in_2')
// (2, 8, 'sp4_h_r_18')
// (3, 7, 'neigh_op_tnr_5')
// (3, 8, 'neigh_op_rgt_5')
// (3, 8, 'sp4_h_r_31')
// (3, 9, 'neigh_op_bnr_5')
// (4, 7, 'neigh_op_top_5')
// (4, 8, 'local_g1_5')
// (4, 8, 'lutff_5/out')
// (4, 8, 'lutff_7/in_1')
// (4, 8, 'sp4_h_r_42')
// (4, 9, 'neigh_op_bot_5')
// (5, 7, 'neigh_op_tnl_5')
// (5, 8, 'neigh_op_lft_5')
// (5, 8, 'sp4_h_l_42')
// (5, 9, 'neigh_op_bnl_5')

reg n75 = 0;
// (1, 8, 'sp4_h_r_9')
// (2, 8, 'local_g1_4')
// (2, 8, 'lutff_7/in_2')
// (2, 8, 'sp4_h_r_20')
// (3, 7, 'neigh_op_tnr_6')
// (3, 8, 'neigh_op_rgt_6')
// (3, 8, 'sp4_h_r_33')
// (3, 9, 'neigh_op_bnr_6')
// (4, 7, 'neigh_op_top_6')
// (4, 8, 'local_g0_6')
// (4, 8, 'lutff_5/in_1')
// (4, 8, 'lutff_6/out')
// (4, 8, 'sp4_h_r_44')
// (4, 9, 'neigh_op_bot_6')
// (5, 7, 'neigh_op_tnl_6')
// (5, 8, 'neigh_op_lft_6')
// (5, 8, 'sp4_h_l_44')
// (5, 9, 'neigh_op_bnl_6')

reg n76 = 0;
// (1, 9, 'neigh_op_tnr_1')
// (1, 10, 'neigh_op_rgt_1')
// (1, 11, 'neigh_op_bnr_1')
// (2, 9, 'neigh_op_top_1')
// (2, 10, 'local_g0_1')
// (2, 10, 'lutff_1/out')
// (2, 10, 'lutff_3/in_0')
// (2, 11, 'neigh_op_bot_1')
// (3, 9, 'neigh_op_tnl_1')
// (3, 10, 'neigh_op_lft_1')
// (3, 11, 'neigh_op_bnl_1')

reg n77 = 0;
// (1, 9, 'sp4_h_r_3')
// (2, 9, 'local_g0_6')
// (2, 9, 'lutff_2/in_0')
// (2, 9, 'sp4_h_r_14')
// (3, 7, 'neigh_op_tnr_3')
// (3, 8, 'neigh_op_rgt_3')
// (3, 9, 'neigh_op_bnr_3')
// (3, 9, 'sp4_h_r_27')
// (4, 6, 'sp4_r_v_b_47')
// (4, 7, 'neigh_op_top_3')
// (4, 7, 'sp4_r_v_b_34')
// (4, 8, 'local_g0_3')
// (4, 8, 'lutff_2/in_1')
// (4, 8, 'lutff_3/out')
// (4, 8, 'sp4_r_v_b_23')
// (4, 9, 'neigh_op_bot_3')
// (4, 9, 'sp4_h_r_38')
// (4, 9, 'sp4_r_v_b_10')
// (5, 5, 'sp4_v_t_47')
// (5, 6, 'sp4_v_b_47')
// (5, 7, 'neigh_op_tnl_3')
// (5, 7, 'sp4_v_b_34')
// (5, 8, 'neigh_op_lft_3')
// (5, 8, 'sp4_v_b_23')
// (5, 9, 'neigh_op_bnl_3')
// (5, 9, 'sp4_h_l_38')
// (5, 9, 'sp4_v_b_10')

wire n78;
// (1, 10, 'local_g0_1')
// (1, 10, 'lutff_5/in_0')
// (1, 10, 'sp4_h_r_9')
// (2, 10, 'sp4_h_r_20')
// (3, 10, 'sp4_h_r_33')
// (4, 7, 'sp4_r_v_b_44')
// (4, 8, 'neigh_op_tnr_2')
// (4, 8, 'sp4_r_v_b_33')
// (4, 9, 'neigh_op_rgt_2')
// (4, 9, 'sp4_r_v_b_20')
// (4, 10, 'neigh_op_bnr_2')
// (4, 10, 'sp4_h_r_44')
// (4, 10, 'sp4_r_v_b_9')
// (5, 6, 'sp4_v_t_44')
// (5, 7, 'sp4_v_b_44')
// (5, 8, 'neigh_op_top_2')
// (5, 8, 'sp4_v_b_33')
// (5, 9, 'local_g1_2')
// (5, 9, 'lutff_2/out')
// (5, 9, 'lutff_3/in_2')
// (5, 9, 'sp4_v_b_20')
// (5, 10, 'local_g0_1')
// (5, 10, 'lutff_1/in_2')
// (5, 10, 'neigh_op_bot_2')
// (5, 10, 'sp4_h_l_44')
// (5, 10, 'sp4_v_b_9')
// (6, 8, 'neigh_op_tnl_2')
// (6, 9, 'neigh_op_lft_2')
// (6, 10, 'neigh_op_bnl_2')

reg n79 = 0;
// (1, 10, 'sp12_h_r_0')
// (2, 10, 'sp12_h_r_3')
// (3, 10, 'sp12_h_r_4')
// (4, 10, 'sp12_h_r_7')
// (5, 10, 'local_g0_0')
// (5, 10, 'lutff_4/in_0')
// (5, 10, 'sp12_h_r_8')
// (6, 9, 'neigh_op_tnr_2')
// (6, 10, 'neigh_op_rgt_2')
// (6, 10, 'sp12_h_r_11')
// (6, 11, 'neigh_op_bnr_2')
// (7, 9, 'neigh_op_top_2')
// (7, 10, 'lutff_2/out')
// (7, 10, 'sp12_h_r_12')
// (7, 11, 'neigh_op_bot_2')
// (8, 9, 'neigh_op_tnl_2')
// (8, 10, 'neigh_op_lft_2')
// (8, 10, 'sp12_h_r_15')
// (8, 11, 'neigh_op_bnl_2')
// (9, 10, 'sp12_h_r_16')
// (10, 10, 'sp12_h_r_19')
// (11, 10, 'sp12_h_r_20')
// (12, 10, 'sp12_h_r_23')
// (13, 10, 'span12_horz_23')

reg n80 = 0;
// (1, 11, 'neigh_op_tnr_0')
// (1, 12, 'neigh_op_rgt_0')
// (1, 13, 'neigh_op_bnr_0')
// (2, 11, 'neigh_op_top_0')
// (2, 12, 'local_g1_0')
// (2, 12, 'lutff_0/out')
// (2, 12, 'lutff_5/in_0')
// (2, 13, 'neigh_op_bot_0')
// (3, 11, 'neigh_op_tnl_0')
// (3, 12, 'neigh_op_lft_0')
// (3, 13, 'neigh_op_bnl_0')

reg n81 = 0;
// (1, 11, 'neigh_op_tnr_5')
// (1, 12, 'neigh_op_rgt_5')
// (1, 13, 'neigh_op_bnr_5')
// (2, 11, 'neigh_op_top_5')
// (2, 12, 'local_g1_5')
// (2, 12, 'lutff_2/in_0')
// (2, 12, 'lutff_5/out')
// (2, 13, 'neigh_op_bot_5')
// (3, 11, 'neigh_op_tnl_5')
// (3, 12, 'neigh_op_lft_5')
// (3, 13, 'neigh_op_bnl_5')

reg n82 = 0;
// (1, 12, 'sp4_h_r_0')
// (2, 12, 'local_g0_5')
// (2, 12, 'lutff_0/in_1')
// (2, 12, 'sp4_h_r_13')
// (3, 10, 'neigh_op_tnr_6')
// (3, 11, 'neigh_op_rgt_6')
// (3, 12, 'neigh_op_bnr_6')
// (3, 12, 'sp4_h_r_24')
// (4, 9, 'sp4_r_v_b_37')
// (4, 10, 'neigh_op_top_6')
// (4, 10, 'sp4_r_v_b_24')
// (4, 11, 'local_g1_6')
// (4, 11, 'lutff_0/in_1')
// (4, 11, 'lutff_6/out')
// (4, 11, 'sp4_r_v_b_13')
// (4, 12, 'neigh_op_bot_6')
// (4, 12, 'sp4_h_r_37')
// (4, 12, 'sp4_r_v_b_0')
// (5, 8, 'sp4_v_t_37')
// (5, 9, 'sp4_v_b_37')
// (5, 10, 'neigh_op_tnl_6')
// (5, 10, 'sp4_v_b_24')
// (5, 11, 'neigh_op_lft_6')
// (5, 11, 'sp4_v_b_13')
// (5, 12, 'neigh_op_bnl_6')
// (5, 12, 'sp4_h_l_37')
// (5, 12, 'sp4_v_b_0')

reg n83 = 0;
// (1, 13, 'neigh_op_tnr_2')
// (1, 14, 'neigh_op_rgt_2')
// (1, 15, 'neigh_op_bnr_2')
// (2, 13, 'neigh_op_top_2')
// (2, 14, 'local_g0_2')
// (2, 14, 'lutff_2/out')
// (2, 14, 'lutff_4/in_0')
// (2, 15, 'neigh_op_bot_2')
// (3, 13, 'neigh_op_tnl_2')
// (3, 14, 'neigh_op_lft_2')
// (3, 15, 'neigh_op_bnl_2')

wire n84;
// (2, 2, 'sp12_h_r_0')
// (3, 2, 'sp12_h_r_3')
// (4, 2, 'sp12_h_r_4')
// (5, 2, 'sp12_h_r_7')
// (6, 2, 'local_g0_0')
// (6, 2, 'local_g1_0')
// (6, 2, 'lutff_1/in_1')
// (6, 2, 'lutff_3/in_2')
// (6, 2, 'lutff_4/in_3')
// (6, 2, 'lutff_6/in_0')
// (6, 2, 'sp12_h_r_8')
// (7, 1, 'local_g2_2')
// (7, 1, 'local_g3_2')
// (7, 1, 'lutff_2/in_0')
// (7, 1, 'lutff_4/in_1')
// (7, 1, 'lutff_5/in_2')
// (7, 1, 'neigh_op_tnr_2')
// (7, 2, 'local_g2_2')
// (7, 2, 'lutff_0/in_0')
// (7, 2, 'neigh_op_rgt_2')
// (7, 2, 'sp12_h_r_11')
// (7, 3, 'neigh_op_bnr_2')
// (8, 1, 'neigh_op_top_2')
// (8, 2, 'lutff_2/out')
// (8, 2, 'sp12_h_r_12')
// (8, 3, 'neigh_op_bot_2')
// (9, 1, 'neigh_op_tnl_2')
// (9, 2, 'neigh_op_lft_2')
// (9, 2, 'sp12_h_r_15')
// (9, 3, 'neigh_op_bnl_2')
// (10, 2, 'sp12_h_r_16')
// (11, 2, 'sp12_h_r_19')
// (12, 2, 'sp12_h_r_20')
// (13, 2, 'span12_horz_20')

wire n85;
// (2, 3, 'lutff_1/cout')
// (2, 3, 'lutff_2/in_3')

wire n86;
// (2, 3, 'lutff_2/cout')
// (2, 3, 'lutff_3/in_3')

wire n87;
// (2, 3, 'lutff_3/cout')
// (2, 3, 'lutff_4/in_3')

wire n88;
// (2, 3, 'lutff_4/cout')
// (2, 3, 'lutff_5/in_3')

wire n89;
// (2, 3, 'lutff_5/cout')
// (2, 3, 'lutff_6/in_3')

wire n90;
// (2, 3, 'lutff_6/cout')
// (2, 3, 'lutff_7/in_3')

wire n91;
// (2, 3, 'sp12_h_r_0')
// (3, 3, 'sp12_h_r_3')
// (4, 3, 'sp12_h_r_4')
// (5, 2, 'sp4_h_r_0')
// (5, 3, 'sp12_h_r_7')
// (6, 2, 'local_g0_5')
// (6, 2, 'lutff_0/in_1')
// (6, 2, 'sp4_h_r_13')
// (6, 3, 'local_g1_0')
// (6, 3, 'lutff_6/in_3')
// (6, 3, 'sp12_h_r_8')
// (7, 2, 'neigh_op_tnr_2')
// (7, 2, 'sp4_h_r_24')
// (7, 3, 'neigh_op_rgt_2')
// (7, 3, 'sp12_h_r_11')
// (7, 4, 'neigh_op_bnr_2')
// (8, 2, 'local_g0_2')
// (8, 2, 'local_g1_2')
// (8, 2, 'lutff_1/in_3')
// (8, 2, 'lutff_7/in_2')
// (8, 2, 'neigh_op_top_2')
// (8, 2, 'sp4_h_r_37')
// (8, 3, 'local_g1_2')
// (8, 3, 'lutff_2/out')
// (8, 3, 'lutff_6/in_1')
// (8, 3, 'sp12_h_r_12')
// (8, 3, 'sp4_r_v_b_37')
// (8, 4, 'neigh_op_bot_2')
// (8, 4, 'sp4_r_v_b_24')
// (8, 5, 'sp4_r_v_b_13')
// (8, 6, 'sp4_r_v_b_0')
// (9, 2, 'neigh_op_tnl_2')
// (9, 2, 'sp4_h_l_37')
// (9, 2, 'sp4_v_t_37')
// (9, 3, 'neigh_op_lft_2')
// (9, 3, 'sp12_h_r_15')
// (9, 3, 'sp4_v_b_37')
// (9, 4, 'neigh_op_bnl_2')
// (9, 4, 'sp4_v_b_24')
// (9, 5, 'sp4_v_b_13')
// (9, 6, 'sp4_v_b_0')
// (10, 3, 'sp12_h_r_16')
// (11, 3, 'sp12_h_r_19')
// (12, 3, 'sp12_h_r_20')
// (13, 3, 'span12_horz_20')

wire n92;
// (2, 4, 'sp12_h_r_1')
// (3, 1, 'sp4_r_v_b_39')
// (3, 2, 'sp4_r_v_b_26')
// (3, 3, 'sp4_r_v_b_15')
// (3, 4, 'sp12_h_r_2')
// (3, 4, 'sp4_r_v_b_2')
// (4, 0, 'span4_vert_39')
// (4, 1, 'sp4_v_b_39')
// (4, 2, 'sp4_v_b_26')
// (4, 3, 'local_g0_7')
// (4, 3, 'lutff_7/in_0')
// (4, 3, 'sp4_v_b_15')
// (4, 4, 'sp12_h_r_5')
// (4, 4, 'sp4_h_r_2')
// (4, 4, 'sp4_v_b_2')
// (5, 1, 'sp4_r_v_b_41')
// (5, 1, 'sp4_r_v_b_44')
// (5, 2, 'sp4_r_v_b_28')
// (5, 2, 'sp4_r_v_b_33')
// (5, 3, 'local_g3_1')
// (5, 3, 'local_g3_4')
// (5, 3, 'lutff_2/in_0')
// (5, 3, 'lutff_4/in_3')
// (5, 3, 'lutff_6/in_3')
// (5, 3, 'sp4_r_v_b_17')
// (5, 3, 'sp4_r_v_b_20')
// (5, 4, 'sp12_h_r_6')
// (5, 4, 'sp4_h_r_15')
// (5, 4, 'sp4_r_v_b_4')
// (5, 4, 'sp4_r_v_b_9')
// (6, 0, 'span4_vert_41')
// (6, 0, 'span4_vert_44')
// (6, 1, 'sp4_v_b_41')
// (6, 1, 'sp4_v_b_44')
// (6, 2, 'sp4_v_b_28')
// (6, 2, 'sp4_v_b_33')
// (6, 3, 'local_g1_4')
// (6, 3, 'lutff_0/in_3')
// (6, 3, 'sp4_v_b_17')
// (6, 3, 'sp4_v_b_20')
// (6, 4, 'sp12_h_r_9')
// (6, 4, 'sp4_h_r_26')
// (6, 4, 'sp4_h_r_4')
// (6, 4, 'sp4_v_b_4')
// (6, 4, 'sp4_v_b_9')
// (7, 1, 'sp4_r_v_b_45')
// (7, 2, 'sp4_r_v_b_32')
// (7, 3, 'local_g3_5')
// (7, 3, 'lutff_0/in_0')
// (7, 3, 'lutff_7/in_3')
// (7, 3, 'sp4_r_v_b_21')
// (7, 4, 'local_g0_2')
// (7, 4, 'lutff_0/in_0')
// (7, 4, 'sp12_h_r_10')
// (7, 4, 'sp4_h_r_17')
// (7, 4, 'sp4_h_r_39')
// (7, 4, 'sp4_r_v_b_8')
// (8, 0, 'span4_vert_45')
// (8, 1, 'sp4_v_b_45')
// (8, 2, 'sp4_v_b_32')
// (8, 3, 'sp4_v_b_21')
// (8, 4, 'sp12_h_r_13')
// (8, 4, 'sp4_h_l_39')
// (8, 4, 'sp4_h_r_28')
// (8, 4, 'sp4_v_b_8')
// (9, 4, 'sp12_h_r_14')
// (9, 4, 'sp4_h_r_41')
// (10, 3, 'neigh_op_tnr_5')
// (10, 4, 'neigh_op_rgt_5')
// (10, 4, 'sp12_h_r_17')
// (10, 4, 'sp4_h_l_41')
// (10, 5, 'neigh_op_bnr_5')
// (11, 3, 'local_g0_5')
// (11, 3, 'lutff_7/in_2')
// (11, 3, 'neigh_op_top_5')
// (11, 4, 'lutff_5/out')
// (11, 4, 'sp12_h_r_18')
// (11, 5, 'neigh_op_bot_5')
// (12, 3, 'neigh_op_tnl_5')
// (12, 4, 'neigh_op_lft_5')
// (12, 4, 'sp12_h_r_21')
// (12, 5, 'neigh_op_bnl_5')
// (13, 4, 'span12_horz_21')

wire n93;
// (2, 5, 'sp12_h_r_1')
// (3, 5, 'sp12_h_r_2')
// (4, 5, 'sp12_h_r_5')
// (5, 5, 'sp12_h_r_6')
// (6, 4, 'neigh_op_tnr_1')
// (6, 5, 'neigh_op_rgt_1')
// (6, 5, 'sp12_h_r_9')
// (6, 6, 'neigh_op_bnr_1')
// (7, 4, 'neigh_op_top_1')
// (7, 5, 'local_g1_2')
// (7, 5, 'lutff_1/out')
// (7, 5, 'lutff_2/in_3')
// (7, 5, 'sp12_h_r_10')
// (7, 6, 'neigh_op_bot_1')
// (8, 4, 'neigh_op_tnl_1')
// (8, 5, 'neigh_op_lft_1')
// (8, 5, 'sp12_h_r_13')
// (8, 6, 'neigh_op_bnl_1')
// (9, 5, 'sp12_h_r_14')
// (10, 5, 'sp12_h_r_17')
// (11, 5, 'sp12_h_r_18')
// (12, 5, 'sp12_h_r_21')
// (13, 5, 'span12_horz_21')

wire n94;
// (2, 6, 'sp4_h_r_8')
// (3, 6, 'sp4_h_r_21')
// (4, 6, 'sp4_h_r_32')
// (5, 3, 'neigh_op_tnr_0')
// (5, 3, 'sp4_r_v_b_45')
// (5, 4, 'neigh_op_rgt_0')
// (5, 4, 'sp4_r_v_b_32')
// (5, 5, 'neigh_op_bnr_0')
// (5, 5, 'sp4_r_v_b_21')
// (5, 6, 'local_g2_0')
// (5, 6, 'local_g2_5')
// (5, 6, 'lutff_1/in_2')
// (5, 6, 'lutff_2/in_2')
// (5, 6, 'lutff_4/in_2')
// (5, 6, 'lutff_7/in_2')
// (5, 6, 'sp4_h_r_45')
// (5, 6, 'sp4_r_v_b_8')
// (6, 2, 'sp4_v_t_45')
// (6, 3, 'neigh_op_top_0')
// (6, 3, 'sp4_v_b_45')
// (6, 4, 'lutff_0/out')
// (6, 4, 'sp4_v_b_32')
// (6, 5, 'neigh_op_bot_0')
// (6, 5, 'sp4_v_b_21')
// (6, 6, 'sp4_h_l_45')
// (6, 6, 'sp4_v_b_8')
// (7, 3, 'neigh_op_tnl_0')
// (7, 4, 'neigh_op_lft_0')
// (7, 5, 'neigh_op_bnl_0')

reg n95 = 0;
// (2, 7, 'sp12_h_r_0')
// (3, 6, 'neigh_op_tnr_6')
// (3, 7, 'neigh_op_rgt_6')
// (3, 7, 'sp12_h_r_3')
// (3, 8, 'neigh_op_bnr_6')
// (4, 6, 'neigh_op_top_6')
// (4, 7, 'lutff_6/out')
// (4, 7, 'sp12_h_r_4')
// (4, 8, 'neigh_op_bot_6')
// (5, 6, 'neigh_op_tnl_6')
// (5, 7, 'neigh_op_lft_6')
// (5, 7, 'sp12_h_r_7')
// (5, 7, 'sp4_h_r_5')
// (5, 8, 'neigh_op_bnl_6')
// (6, 7, 'local_g1_0')
// (6, 7, 'lutff_1/in_0')
// (6, 7, 'sp12_h_r_8')
// (6, 7, 'sp4_h_r_16')
// (7, 7, 'local_g2_5')
// (7, 7, 'lutff_6/in_1')
// (7, 7, 'sp12_h_r_11')
// (7, 7, 'sp4_h_r_29')
// (8, 7, 'sp12_h_r_12')
// (8, 7, 'sp4_h_r_40')
// (9, 7, 'sp12_h_r_15')
// (9, 7, 'sp4_h_l_40')
// (10, 7, 'sp12_h_r_16')
// (11, 7, 'sp12_h_r_19')
// (12, 7, 'sp12_h_r_20')
// (13, 7, 'span12_horz_20')

reg n96 = 0;
// (2, 10, 'sp4_h_r_8')
// (3, 10, 'sp4_h_r_21')
// (4, 10, 'sp4_h_r_32')
// (5, 10, 'sp4_h_r_45')
// (5, 11, 'sp4_r_v_b_36')
// (5, 11, 'sp4_r_v_b_39')
// (5, 12, 'local_g0_1')
// (5, 12, 'local_g0_2')
// (5, 12, 'lutff_4/in_2')
// (5, 12, 'lutff_5/in_2')
// (5, 12, 'sp4_r_v_b_25')
// (5, 12, 'sp4_r_v_b_26')
// (5, 13, 'sp4_r_v_b_12')
// (5, 13, 'sp4_r_v_b_15')
// (5, 14, 'sp4_r_v_b_1')
// (5, 14, 'sp4_r_v_b_2')
// (6, 10, 'sp4_h_l_45')
// (6, 10, 'sp4_h_r_8')
// (6, 10, 'sp4_v_t_36')
// (6, 10, 'sp4_v_t_39')
// (6, 11, 'sp4_v_b_36')
// (6, 11, 'sp4_v_b_39')
// (6, 12, 'sp4_v_b_25')
// (6, 12, 'sp4_v_b_26')
// (6, 13, 'sp4_v_b_12')
// (6, 13, 'sp4_v_b_15')
// (6, 14, 'sp4_v_b_1')
// (6, 14, 'sp4_v_b_2')
// (7, 10, 'sp4_h_r_21')
// (8, 6, 'neigh_op_tnr_6')
// (8, 7, 'neigh_op_rgt_6')
// (8, 8, 'neigh_op_bnr_6')
// (8, 10, 'sp4_h_r_32')
// (9, 1, 'sp12_v_t_23')
// (9, 2, 'sp12_v_b_23')
// (9, 3, 'sp12_v_b_20')
// (9, 4, 'sp12_v_b_19')
// (9, 5, 'sp12_v_b_16')
// (9, 6, 'neigh_op_top_6')
// (9, 6, 'sp12_v_b_15')
// (9, 7, 'lutff_6/out')
// (9, 7, 'sp12_v_b_12')
// (9, 7, 'sp4_r_v_b_45')
// (9, 8, 'neigh_op_bot_6')
// (9, 8, 'sp12_v_b_11')
// (9, 8, 'sp4_r_v_b_32')
// (9, 9, 'sp12_v_b_8')
// (9, 9, 'sp4_r_v_b_21')
// (9, 10, 'sp12_v_b_7')
// (9, 10, 'sp4_h_r_45')
// (9, 10, 'sp4_r_v_b_8')
// (9, 11, 'sp12_v_b_4')
// (9, 12, 'local_g3_3')
// (9, 12, 'lutff_4/in_0')
// (9, 12, 'sp12_v_b_3')
// (9, 13, 'sp12_v_b_0')
// (10, 6, 'neigh_op_tnl_6')
// (10, 6, 'sp4_h_r_1')
// (10, 6, 'sp4_v_t_45')
// (10, 7, 'neigh_op_lft_6')
// (10, 7, 'sp4_v_b_45')
// (10, 8, 'neigh_op_bnl_6')
// (10, 8, 'sp4_v_b_32')
// (10, 9, 'sp4_v_b_21')
// (10, 10, 'sp4_h_l_45')
// (10, 10, 'sp4_v_b_8')
// (11, 6, 'local_g0_4')
// (11, 6, 'lutff_6/in_0')
// (11, 6, 'sp4_h_r_12')
// (12, 6, 'sp4_h_r_25')
// (13, 6, 'span4_horz_25')

wire n97;
// (2, 11, 'sp12_h_r_0')
// (3, 11, 'sp12_h_r_3')
// (4, 11, 'sp12_h_r_4')
// (5, 10, 'neigh_op_tnr_0')
// (5, 11, 'neigh_op_rgt_0')
// (5, 11, 'sp12_h_r_7')
// (5, 12, 'neigh_op_bnr_0')
// (6, 10, 'neigh_op_top_0')
// (6, 11, 'lutff_0/out')
// (6, 11, 'sp12_h_r_8')
// (6, 12, 'neigh_op_bot_0')
// (7, 10, 'neigh_op_tnl_0')
// (7, 11, 'local_g1_0')
// (7, 11, 'lutff_2/in_1')
// (7, 11, 'neigh_op_lft_0')
// (7, 11, 'sp12_h_r_11')
// (7, 12, 'neigh_op_bnl_0')
// (8, 11, 'local_g0_4')
// (8, 11, 'lutff_3/in_1')
// (8, 11, 'sp12_h_r_12')
// (9, 11, 'sp12_h_r_15')
// (10, 11, 'sp12_h_r_16')
// (11, 11, 'sp12_h_r_19')
// (12, 11, 'sp12_h_r_20')
// (13, 11, 'span12_horz_20')

reg n98 = 0;
// (2, 12, 'local_g0_2')
// (2, 12, 'lutff_0/in_0')
// (2, 12, 'sp4_h_r_10')
// (3, 11, 'neigh_op_tnr_1')
// (3, 12, 'neigh_op_rgt_1')
// (3, 12, 'sp4_h_r_23')
// (3, 13, 'neigh_op_bnr_1')
// (4, 11, 'local_g0_1')
// (4, 11, 'lutff_1/in_0')
// (4, 11, 'lutff_3/in_0')
// (4, 11, 'neigh_op_top_1')
// (4, 12, 'local_g1_1')
// (4, 12, 'lutff_1/out')
// (4, 12, 'lutff_6/in_0')
// (4, 12, 'sp4_h_r_34')
// (4, 13, 'neigh_op_bot_1')
// (5, 11, 'neigh_op_tnl_1')
// (5, 12, 'neigh_op_lft_1')
// (5, 12, 'sp4_h_r_47')
// (5, 13, 'neigh_op_bnl_1')
// (6, 12, 'sp4_h_l_47')

reg n99 = 0;
// (2, 13, 'local_g0_2')
// (2, 13, 'lutff_4/in_0')
// (2, 13, 'sp4_h_r_10')
// (3, 12, 'neigh_op_tnr_1')
// (3, 13, 'neigh_op_rgt_1')
// (3, 13, 'sp4_h_r_23')
// (3, 14, 'neigh_op_bnr_1')
// (4, 12, 'neigh_op_top_1')
// (4, 13, 'lutff_1/out')
// (4, 13, 'sp4_h_r_34')
// (4, 14, 'neigh_op_bot_1')
// (5, 12, 'neigh_op_tnl_1')
// (5, 13, 'neigh_op_lft_1')
// (5, 13, 'sp4_h_r_47')
// (5, 14, 'neigh_op_bnl_1')
// (6, 13, 'sp4_h_l_47')

reg n100 = 0;
// (2, 13, 'sp12_h_r_0')
// (3, 13, 'sp12_h_r_3')
// (4, 13, 'sp12_h_r_4')
// (5, 13, 'sp12_h_r_7')
// (6, 13, 'sp12_h_r_8')
// (7, 12, 'neigh_op_tnr_2')
// (7, 13, 'neigh_op_rgt_2')
// (7, 13, 'sp12_h_r_11')
// (7, 14, 'neigh_op_bnr_2')
// (8, 12, 'neigh_op_top_2')
// (8, 13, 'lutff_2/out')
// (8, 13, 'sp12_h_r_12')
// (8, 14, 'neigh_op_bot_2')
// (9, 12, 'neigh_op_tnl_2')
// (9, 13, 'neigh_op_lft_2')
// (9, 13, 'sp12_h_r_15')
// (9, 14, 'neigh_op_bnl_2')
// (10, 13, 'sp12_h_r_16')
// (11, 13, 'local_g1_3')
// (11, 13, 'lutff_4/in_0')
// (11, 13, 'sp12_h_r_19')
// (12, 13, 'sp12_h_r_20')
// (13, 13, 'span12_horz_20')

reg n101 = 0;
// (3, 1, 'sp4_r_v_b_47')
// (3, 2, 'sp4_r_v_b_34')
// (3, 3, 'neigh_op_tnr_5')
// (3, 3, 'sp4_r_v_b_23')
// (3, 4, 'neigh_op_rgt_5')
// (3, 4, 'sp4_r_v_b_10')
// (3, 5, 'neigh_op_bnr_5')
// (4, 0, 'span4_vert_47')
// (4, 1, 'sp4_v_b_47')
// (4, 2, 'sp4_v_b_34')
// (4, 3, 'local_g1_7')
// (4, 3, 'lutff_7/in_3')
// (4, 3, 'neigh_op_top_5')
// (4, 3, 'sp4_v_b_23')
// (4, 4, 'lutff_5/out')
// (4, 4, 'sp4_v_b_10')
// (4, 5, 'neigh_op_bot_5')
// (5, 3, 'neigh_op_tnl_5')
// (5, 4, 'neigh_op_lft_5')
// (5, 5, 'neigh_op_bnl_5')

wire n102;
// (3, 2, 'neigh_op_tnr_1')
// (3, 3, 'neigh_op_rgt_1')
// (3, 4, 'neigh_op_bnr_1')
// (4, 2, 'neigh_op_top_1')
// (4, 3, 'local_g0_1')
// (4, 3, 'lutff_1/out')
// (4, 3, 'lutff_7/in_2')
// (4, 4, 'neigh_op_bot_1')
// (5, 2, 'neigh_op_tnl_1')
// (5, 3, 'neigh_op_lft_1')
// (5, 4, 'neigh_op_bnl_1')

wire n103;
// (3, 2, 'neigh_op_tnr_2')
// (3, 3, 'neigh_op_rgt_2')
// (3, 4, 'neigh_op_bnr_2')
// (4, 2, 'neigh_op_top_2')
// (4, 3, 'lutff_2/out')
// (4, 4, 'neigh_op_bot_2')
// (5, 2, 'neigh_op_tnl_2')
// (5, 3, 'local_g0_2')
// (5, 3, 'lutff_4/in_2')
// (5, 3, 'neigh_op_lft_2')
// (5, 4, 'neigh_op_bnl_2')

wire n104;
// (3, 2, 'neigh_op_tnr_5')
// (3, 3, 'neigh_op_rgt_5')
// (3, 4, 'neigh_op_bnr_5')
// (4, 2, 'neigh_op_top_5')
// (4, 3, 'local_g1_5')
// (4, 3, 'local_g2_5')
// (4, 3, 'lutff_1/in_0')
// (4, 3, 'lutff_2/in_2')
// (4, 3, 'lutff_5/out')
// (4, 4, 'neigh_op_bot_5')
// (5, 2, 'neigh_op_tnl_5')
// (5, 3, 'neigh_op_lft_5')
// (5, 4, 'neigh_op_bnl_5')

wire n105;
// (3, 2, 'sp4_h_r_2')
// (4, 1, 'neigh_op_tnr_5')
// (4, 2, 'neigh_op_rgt_5')
// (4, 2, 'sp4_h_r_15')
// (4, 3, 'neigh_op_bnr_5')
// (5, 1, 'neigh_op_top_5')
// (5, 2, 'lutff_5/out')
// (5, 2, 'sp4_h_r_26')
// (5, 3, 'neigh_op_bot_5')
// (6, 1, 'neigh_op_tnl_5')
// (6, 1, 'sp4_r_v_b_15')
// (6, 2, 'neigh_op_lft_5')
// (6, 2, 'sp4_h_r_39')
// (6, 2, 'sp4_r_v_b_2')
// (6, 3, 'neigh_op_bnl_5')
// (6, 3, 'sp4_r_v_b_40')
// (6, 4, 'sp4_r_v_b_29')
// (6, 5, 'sp4_r_v_b_16')
// (6, 6, 'sp4_r_v_b_5')
// (7, 0, 'span4_vert_15')
// (7, 1, 'sp4_v_b_15')
// (7, 2, 'sp4_h_l_39')
// (7, 2, 'sp4_v_b_2')
// (7, 2, 'sp4_v_t_40')
// (7, 3, 'local_g2_0')
// (7, 3, 'lutff_0/in_2')
// (7, 3, 'sp4_v_b_40')
// (7, 4, 'sp4_v_b_29')
// (7, 5, 'sp4_v_b_16')
// (7, 6, 'sp4_v_b_5')

reg n106 = 0;
// (3, 3, 'neigh_op_tnr_0')
// (3, 4, 'neigh_op_rgt_0')
// (3, 5, 'neigh_op_bnr_0')
// (4, 3, 'neigh_op_top_0')
// (4, 4, 'local_g1_0')
// (4, 4, 'lutff_0/out')
// (4, 4, 'lutff_5/in_0')
// (4, 5, 'neigh_op_bot_0')
// (5, 3, 'neigh_op_tnl_0')
// (5, 4, 'neigh_op_lft_0')
// (5, 5, 'neigh_op_bnl_0')

reg n107 = 0;
// (3, 3, 'neigh_op_tnr_7')
// (3, 4, 'neigh_op_rgt_7')
// (3, 5, 'neigh_op_bnr_7')
// (4, 3, 'neigh_op_top_7')
// (4, 4, 'local_g1_7')
// (4, 4, 'lutff_0/in_0')
// (4, 4, 'lutff_7/out')
// (4, 5, 'neigh_op_bot_7')
// (5, 3, 'neigh_op_tnl_7')
// (5, 4, 'neigh_op_lft_7')
// (5, 5, 'neigh_op_bnl_7')

wire n108;
// (3, 3, 'sp12_h_r_1')
// (4, 3, 'sp12_h_r_2')
// (5, 3, 'sp12_h_r_5')
// (6, 3, 'sp12_h_r_6')
// (7, 2, 'local_g2_1')
// (7, 2, 'local_g3_1')
// (7, 2, 'lutff_1/in_0')
// (7, 2, 'lutff_2/in_0')
// (7, 2, 'neigh_op_tnr_1')
// (7, 3, 'local_g1_1')
// (7, 3, 'lutff_3/in_3')
// (7, 3, 'lutff_5/in_3')
// (7, 3, 'neigh_op_rgt_1')
// (7, 3, 'sp12_h_r_9')
// (7, 4, 'neigh_op_bnr_1')
// (8, 2, 'local_g1_1')
// (8, 2, 'lutff_2/in_0')
// (8, 2, 'neigh_op_top_1')
// (8, 3, 'lutff_1/out')
// (8, 3, 'sp12_h_r_10')
// (8, 4, 'neigh_op_bot_1')
// (9, 2, 'neigh_op_tnl_1')
// (9, 3, 'neigh_op_lft_1')
// (9, 3, 'sp12_h_r_13')
// (9, 4, 'neigh_op_bnl_1')
// (10, 3, 'sp12_h_r_14')
// (11, 3, 'sp12_h_r_17')
// (12, 3, 'sp12_h_r_18')
// (13, 3, 'span12_horz_18')

wire n109;
// (3, 3, 'sp4_h_r_4')
// (4, 3, 'sp4_h_r_17')
// (5, 3, 'sp4_h_r_28')
// (6, 3, 'local_g2_1')
// (6, 3, 'local_g3_1')
// (6, 3, 'lutff_2/in_3')
// (6, 3, 'lutff_7/in_3')
// (6, 3, 'sp4_h_r_41')
// (7, 3, 'sp4_h_l_41')
// (7, 3, 'sp4_h_r_8')
// (8, 3, 'sp4_h_r_21')
// (9, 3, 'sp4_h_r_32')
// (10, 1, 'neigh_op_tnr_7')
// (10, 1, 'sp4_r_v_b_27')
// (10, 2, 'neigh_op_rgt_7')
// (10, 2, 'sp4_r_v_b_14')
// (10, 3, 'neigh_op_bnr_7')
// (10, 3, 'sp4_h_r_45')
// (10, 3, 'sp4_r_v_b_3')
// (11, 0, 'span4_vert_27')
// (11, 1, 'neigh_op_top_7')
// (11, 1, 'sp4_v_b_27')
// (11, 2, 'lutff_7/out')
// (11, 2, 'sp4_v_b_14')
// (11, 3, 'neigh_op_bot_7')
// (11, 3, 'sp4_h_l_45')
// (11, 3, 'sp4_v_b_3')
// (12, 1, 'neigh_op_tnl_7')
// (12, 2, 'neigh_op_lft_7')
// (12, 3, 'neigh_op_bnl_7')

reg n110 = 0;
// (3, 4, 'neigh_op_tnr_0')
// (3, 5, 'neigh_op_rgt_0')
// (3, 6, 'neigh_op_bnr_0')
// (4, 4, 'neigh_op_top_0')
// (4, 5, 'local_g3_0')
// (4, 5, 'lutff_0/out')
// (4, 5, 'lutff_5/in_0')
// (4, 6, 'neigh_op_bot_0')
// (5, 4, 'neigh_op_tnl_0')
// (5, 5, 'neigh_op_lft_0')
// (5, 6, 'neigh_op_bnl_0')

reg \d_out[6] = 0 ;
// (3, 4, 'neigh_op_tnr_3')
// (3, 5, 'neigh_op_rgt_3')
// (3, 6, 'neigh_op_bnr_3')
// (4, 0, 'io_1/D_OUT_0')
// (4, 0, 'io_1/PAD')
// (4, 0, 'local_g1_6')
// (4, 0, 'span12_vert_14')
// (4, 1, 'sp12_v_b_14')
// (4, 2, 'sp12_v_b_13')
// (4, 3, 'sp12_v_b_10')
// (4, 4, 'neigh_op_top_3')
// (4, 4, 'sp12_v_b_9')
// (4, 5, 'lutff_3/out')
// (4, 5, 'sp12_v_b_6')
// (4, 6, 'neigh_op_bot_3')
// (4, 6, 'sp12_v_b_5')
// (4, 7, 'sp12_v_b_2')
// (4, 8, 'sp12_v_b_1')
// (5, 4, 'neigh_op_tnl_3')
// (5, 5, 'neigh_op_lft_3')
// (5, 6, 'neigh_op_bnl_3')

reg n112 = 0;
// (3, 4, 'neigh_op_tnr_4')
// (3, 5, 'neigh_op_rgt_4')
// (3, 6, 'neigh_op_bnr_4')
// (4, 4, 'neigh_op_top_4')
// (4, 5, 'local_g0_4')
// (4, 5, 'lutff_0/in_0')
// (4, 5, 'lutff_4/out')
// (4, 6, 'neigh_op_bot_4')
// (5, 4, 'neigh_op_tnl_4')
// (5, 5, 'neigh_op_lft_4')
// (5, 6, 'neigh_op_bnl_4')

reg n113 = 0;
// (3, 4, 'neigh_op_tnr_5')
// (3, 5, 'neigh_op_rgt_5')
// (3, 6, 'neigh_op_bnr_5')
// (4, 4, 'neigh_op_top_5')
// (4, 5, 'local_g1_5')
// (4, 5, 'lutff_2/in_0')
// (4, 5, 'lutff_5/out')
// (4, 6, 'neigh_op_bot_5')
// (5, 4, 'neigh_op_tnl_5')
// (5, 5, 'neigh_op_lft_5')
// (5, 6, 'neigh_op_bnl_5')

reg n114 = 0;
// (3, 4, 'neigh_op_tnr_7')
// (3, 5, 'neigh_op_rgt_7')
// (3, 6, 'neigh_op_bnr_7')
// (4, 4, 'local_g0_7')
// (4, 4, 'lutff_7/in_0')
// (4, 4, 'neigh_op_top_7')
// (4, 5, 'lutff_7/out')
// (4, 6, 'neigh_op_bot_7')
// (5, 4, 'neigh_op_tnl_7')
// (5, 5, 'neigh_op_lft_7')
// (5, 6, 'neigh_op_bnl_7')

wire n115;
// (3, 4, 'sp12_h_r_0')
// (4, 4, 'sp12_h_r_3')
// (5, 4, 'sp12_h_r_4')
// (6, 4, 'sp12_h_r_7')
// (7, 4, 'sp12_h_r_8')
// (8, 3, 'neigh_op_tnr_2')
// (8, 4, 'neigh_op_rgt_2')
// (8, 4, 'sp12_h_r_11')
// (8, 5, 'neigh_op_bnr_2')
// (9, 3, 'neigh_op_top_2')
// (9, 4, 'lutff_2/out')
// (9, 4, 'sp12_h_r_12')
// (9, 5, 'neigh_op_bot_2')
// (10, 3, 'neigh_op_tnl_2')
// (10, 4, 'neigh_op_lft_2')
// (10, 4, 'sp12_h_r_15')
// (10, 5, 'neigh_op_bnl_2')
// (11, 4, 'local_g1_0')
// (11, 4, 'lutff_1/in_2')
// (11, 4, 'lutff_7/in_2')
// (11, 4, 'sp12_h_r_16')
// (12, 4, 'sp12_h_r_19')
// (13, 4, 'span12_horz_19')

reg n116 = 0;
// (3, 4, 'sp4_r_v_b_43')
// (3, 5, 'sp4_r_v_b_30')
// (3, 6, 'sp4_r_v_b_19')
// (3, 7, 'sp4_r_v_b_6')
// (4, 3, 'sp4_v_t_43')
// (4, 4, 'sp4_v_b_43')
// (4, 5, 'local_g2_6')
// (4, 5, 'lutff_7/in_3')
// (4, 5, 'sp4_v_b_30')
// (4, 6, 'neigh_op_tnr_6')
// (4, 6, 'sp4_v_b_19')
// (4, 7, 'neigh_op_rgt_6')
// (4, 7, 'sp4_h_r_1')
// (4, 7, 'sp4_v_b_6')
// (4, 8, 'neigh_op_bnr_6')
// (5, 6, 'neigh_op_top_6')
// (5, 7, 'lutff_6/out')
// (5, 7, 'sp4_h_r_12')
// (5, 8, 'neigh_op_bot_6')
// (6, 6, 'neigh_op_tnl_6')
// (6, 7, 'neigh_op_lft_6')
// (6, 7, 'sp4_h_r_25')
// (6, 8, 'neigh_op_bnl_6')
// (7, 7, 'sp4_h_r_36')
// (8, 7, 'sp4_h_l_36')

reg \d_out[7] = 0 ;
// (3, 5, 'neigh_op_tnr_0')
// (3, 6, 'neigh_op_rgt_0')
// (3, 7, 'neigh_op_bnr_0')
// (4, 0, 'io_0/D_OUT_0')
// (4, 0, 'io_0/PAD')
// (4, 0, 'local_g1_3')
// (4, 0, 'span12_vert_11')
// (4, 1, 'sp12_v_b_11')
// (4, 2, 'sp12_v_b_8')
// (4, 3, 'sp12_v_b_7')
// (4, 4, 'sp12_v_b_4')
// (4, 5, 'neigh_op_top_0')
// (4, 5, 'sp12_v_b_3')
// (4, 6, 'lutff_0/out')
// (4, 6, 'sp12_v_b_0')
// (4, 7, 'neigh_op_bot_0')
// (5, 5, 'neigh_op_tnl_0')
// (5, 6, 'neigh_op_lft_0')
// (5, 7, 'neigh_op_bnl_0')

reg n118 = 0;
// (3, 5, 'neigh_op_tnr_2')
// (3, 6, 'neigh_op_rgt_2')
// (3, 7, 'neigh_op_bnr_2')
// (4, 5, 'local_g1_2')
// (4, 5, 'lutff_4/in_3')
// (4, 5, 'neigh_op_top_2')
// (4, 6, 'lutff_2/out')
// (4, 7, 'neigh_op_bot_2')
// (5, 5, 'neigh_op_tnl_2')
// (5, 6, 'neigh_op_lft_2')
// (5, 7, 'neigh_op_bnl_2')

reg n119 = 0;
// (3, 5, 'neigh_op_tnr_3')
// (3, 6, 'neigh_op_rgt_3')
// (3, 7, 'neigh_op_bnr_3')
// (4, 5, 'neigh_op_top_3')
// (4, 6, 'local_g0_3')
// (4, 6, 'lutff_3/out')
// (4, 6, 'lutff_7/in_0')
// (4, 7, 'neigh_op_bot_3')
// (5, 5, 'neigh_op_tnl_3')
// (5, 6, 'neigh_op_lft_3')
// (5, 7, 'neigh_op_bnl_3')

reg n120 = 0;
// (3, 5, 'neigh_op_tnr_4')
// (3, 6, 'neigh_op_rgt_4')
// (3, 7, 'neigh_op_bnr_4')
// (4, 5, 'neigh_op_top_4')
// (4, 6, 'lutff_4/out')
// (4, 6, 'sp4_h_r_8')
// (4, 7, 'neigh_op_bot_4')
// (5, 5, 'neigh_op_tnl_4')
// (5, 6, 'neigh_op_lft_4')
// (5, 6, 'sp4_h_r_21')
// (5, 7, 'neigh_op_bnl_4')
// (6, 6, 'sp4_h_r_32')
// (7, 6, 'sp4_h_r_45')
// (7, 7, 'local_g3_5')
// (7, 7, 'lutff_2/in_0')
// (7, 7, 'sp4_r_v_b_45')
// (7, 8, 'sp4_r_v_b_32')
// (7, 9, 'sp4_r_v_b_21')
// (7, 10, 'sp4_r_v_b_8')
// (8, 6, 'sp4_h_l_45')
// (8, 6, 'sp4_v_t_45')
// (8, 7, 'sp4_v_b_45')
// (8, 8, 'sp4_v_b_32')
// (8, 9, 'sp4_v_b_21')
// (8, 10, 'sp4_v_b_8')

reg n121 = 0;
// (3, 6, 'neigh_op_tnr_4')
// (3, 7, 'neigh_op_rgt_4')
// (3, 8, 'neigh_op_bnr_4')
// (4, 6, 'neigh_op_top_4')
// (4, 7, 'local_g0_4')
// (4, 7, 'lutff_4/out')
// (4, 7, 'lutff_6/in_0')
// (4, 8, 'neigh_op_bot_4')
// (5, 6, 'neigh_op_tnl_4')
// (5, 7, 'neigh_op_lft_4')
// (5, 8, 'neigh_op_bnl_4')

wire n122;
// (3, 6, 'sp4_h_r_1')
// (4, 6, 'sp4_h_r_12')
// (5, 4, 'neigh_op_tnr_2')
// (5, 5, 'local_g3_2')
// (5, 5, 'lutff_0/in_1')
// (5, 5, 'neigh_op_rgt_2')
// (5, 6, 'local_g3_1')
// (5, 6, 'lutff_3/in_3')
// (5, 6, 'neigh_op_bnr_2')
// (5, 6, 'sp4_h_r_25')
// (6, 3, 'sp4_r_v_b_45')
// (6, 4, 'neigh_op_top_2')
// (6, 4, 'sp4_r_v_b_32')
// (6, 5, 'lutff_2/out')
// (6, 5, 'sp4_r_v_b_21')
// (6, 6, 'neigh_op_bot_2')
// (6, 6, 'sp4_h_r_36')
// (6, 6, 'sp4_r_v_b_8')
// (7, 2, 'sp4_v_t_45')
// (7, 3, 'sp4_v_b_45')
// (7, 4, 'neigh_op_tnl_2')
// (7, 4, 'sp4_v_b_32')
// (7, 5, 'neigh_op_lft_2')
// (7, 5, 'sp4_v_b_21')
// (7, 6, 'neigh_op_bnl_2')
// (7, 6, 'sp4_h_l_36')
// (7, 6, 'sp4_v_b_8')

wire n123;
// (3, 6, 'sp4_h_r_4')
// (4, 6, 'sp4_h_r_17')
// (5, 4, 'neigh_op_tnr_0')
// (5, 5, 'local_g3_0')
// (5, 5, 'lutff_5/in_0')
// (5, 5, 'neigh_op_rgt_0')
// (5, 6, 'local_g2_4')
// (5, 6, 'lutff_0/in_0')
// (5, 6, 'lutff_3/in_1')
// (5, 6, 'lutff_6/in_0')
// (5, 6, 'neigh_op_bnr_0')
// (5, 6, 'sp4_h_r_28')
// (6, 3, 'sp4_r_v_b_41')
// (6, 4, 'neigh_op_top_0')
// (6, 4, 'sp4_r_v_b_28')
// (6, 5, 'lutff_0/out')
// (6, 5, 'sp4_r_v_b_17')
// (6, 6, 'neigh_op_bot_0')
// (6, 6, 'sp4_h_r_41')
// (6, 6, 'sp4_r_v_b_4')
// (7, 2, 'sp4_v_t_41')
// (7, 3, 'sp4_v_b_41')
// (7, 4, 'neigh_op_tnl_0')
// (7, 4, 'sp4_v_b_28')
// (7, 5, 'neigh_op_lft_0')
// (7, 5, 'sp4_v_b_17')
// (7, 6, 'neigh_op_bnl_0')
// (7, 6, 'sp4_h_l_41')
// (7, 6, 'sp4_v_b_4')

reg n124 = 0;
// (3, 7, 'neigh_op_tnr_4')
// (3, 8, 'neigh_op_rgt_4')
// (3, 9, 'neigh_op_bnr_4')
// (4, 7, 'neigh_op_top_4')
// (4, 7, 'sp4_r_v_b_36')
// (4, 8, 'lutff_4/out')
// (4, 8, 'sp4_r_v_b_25')
// (4, 9, 'local_g2_4')
// (4, 9, 'lutff_1/in_1')
// (4, 9, 'lutff_6/in_2')
// (4, 9, 'neigh_op_bot_4')
// (4, 9, 'sp4_r_v_b_12')
// (4, 10, 'sp4_r_v_b_1')
// (5, 6, 'sp4_v_t_36')
// (5, 7, 'neigh_op_tnl_4')
// (5, 7, 'sp4_v_b_36')
// (5, 8, 'neigh_op_lft_4')
// (5, 8, 'sp4_v_b_25')
// (5, 9, 'neigh_op_bnl_4')
// (5, 9, 'sp4_v_b_12')
// (5, 10, 'sp4_v_b_1')

reg n125 = 0;
// (3, 7, 'neigh_op_tnr_7')
// (3, 8, 'neigh_op_rgt_7')
// (3, 9, 'neigh_op_bnr_7')
// (4, 7, 'neigh_op_top_7')
// (4, 8, 'local_g1_7')
// (4, 8, 'lutff_0/in_2')
// (4, 8, 'lutff_1/in_1')
// (4, 8, 'lutff_7/out')
// (4, 9, 'neigh_op_bot_7')
// (5, 7, 'neigh_op_tnl_7')
// (5, 8, 'neigh_op_lft_7')
// (5, 9, 'neigh_op_bnl_7')

reg n126 = 0;
// (3, 8, 'neigh_op_tnr_0')
// (3, 9, 'neigh_op_rgt_0')
// (3, 10, 'neigh_op_bnr_0')
// (4, 8, 'neigh_op_top_0')
// (4, 9, 'local_g3_0')
// (4, 9, 'lutff_0/out')
// (4, 9, 'lutff_4/in_1')
// (4, 10, 'neigh_op_bot_0')
// (5, 8, 'neigh_op_tnl_0')
// (5, 9, 'neigh_op_lft_0')
// (5, 10, 'neigh_op_bnl_0')

reg n127 = 0;
// (3, 8, 'neigh_op_tnr_1')
// (3, 9, 'neigh_op_rgt_1')
// (3, 10, 'neigh_op_bnr_1')
// (4, 8, 'local_g1_1')
// (4, 8, 'lutff_3/in_1')
// (4, 8, 'neigh_op_top_1')
// (4, 9, 'lutff_1/out')
// (4, 10, 'local_g0_1')
// (4, 10, 'lutff_3/in_2')
// (4, 10, 'neigh_op_bot_1')
// (5, 8, 'neigh_op_tnl_1')
// (5, 9, 'neigh_op_lft_1')
// (5, 10, 'neigh_op_bnl_1')

reg n128 = 0;
// (3, 8, 'neigh_op_tnr_2')
// (3, 9, 'neigh_op_rgt_2')
// (3, 10, 'neigh_op_bnr_2')
// (4, 8, 'neigh_op_top_2')
// (4, 9, 'local_g0_2')
// (4, 9, 'lutff_0/in_2')
// (4, 9, 'lutff_2/out')
// (4, 9, 'lutff_3/in_1')
// (4, 10, 'neigh_op_bot_2')
// (5, 8, 'neigh_op_tnl_2')
// (5, 9, 'neigh_op_lft_2')
// (5, 10, 'neigh_op_bnl_2')

reg n129 = 0;
// (3, 8, 'neigh_op_tnr_3')
// (3, 9, 'neigh_op_rgt_3')
// (3, 10, 'neigh_op_bnr_3')
// (4, 8, 'neigh_op_top_3')
// (4, 9, 'local_g1_3')
// (4, 9, 'lutff_3/out')
// (4, 9, 'lutff_4/in_2')
// (4, 9, 'lutff_5/in_1')
// (4, 10, 'neigh_op_bot_3')
// (5, 8, 'neigh_op_tnl_3')
// (5, 9, 'neigh_op_lft_3')
// (5, 10, 'neigh_op_bnl_3')

reg n130 = 0;
// (3, 8, 'neigh_op_tnr_4')
// (3, 9, 'neigh_op_rgt_4')
// (3, 10, 'neigh_op_bnr_4')
// (4, 8, 'neigh_op_top_4')
// (4, 9, 'lutff_4/out')
// (4, 10, 'local_g1_4')
// (4, 10, 'lutff_2/in_1')
// (4, 10, 'neigh_op_bot_4')
// (5, 8, 'neigh_op_tnl_4')
// (5, 9, 'neigh_op_lft_4')
// (5, 10, 'neigh_op_bnl_4')

reg n131 = 0;
// (3, 8, 'neigh_op_tnr_5')
// (3, 9, 'neigh_op_rgt_5')
// (3, 10, 'neigh_op_bnr_5')
// (4, 8, 'neigh_op_top_5')
// (4, 9, 'local_g0_5')
// (4, 9, 'lutff_5/out')
// (4, 9, 'lutff_7/in_0')
// (4, 10, 'local_g1_5')
// (4, 10, 'lutff_2/in_2')
// (4, 10, 'neigh_op_bot_5')
// (5, 8, 'neigh_op_tnl_5')
// (5, 9, 'neigh_op_lft_5')
// (5, 10, 'neigh_op_bnl_5')

reg n132 = 0;
// (3, 8, 'neigh_op_tnr_6')
// (3, 9, 'neigh_op_rgt_6')
// (3, 10, 'neigh_op_bnr_6')
// (4, 8, 'neigh_op_top_6')
// (4, 9, 'lutff_6/out')
// (4, 10, 'local_g0_6')
// (4, 10, 'lutff_3/in_1')
// (4, 10, 'neigh_op_bot_6')
// (5, 8, 'neigh_op_tnl_6')
// (5, 9, 'neigh_op_lft_6')
// (5, 10, 'neigh_op_bnl_6')

wire n133;
// (3, 8, 'sp4_r_v_b_38')
// (3, 9, 'neigh_op_tnr_7')
// (3, 9, 'sp4_r_v_b_27')
// (3, 10, 'neigh_op_rgt_7')
// (3, 10, 'sp4_r_v_b_14')
// (3, 11, 'neigh_op_bnr_7')
// (3, 11, 'sp4_r_v_b_3')
// (4, 7, 'sp4_h_r_3')
// (4, 7, 'sp4_v_t_38')
// (4, 8, 'sp4_v_b_38')
// (4, 9, 'neigh_op_top_7')
// (4, 9, 'sp4_v_b_27')
// (4, 10, 'lutff_7/out')
// (4, 10, 'sp4_v_b_14')
// (4, 11, 'neigh_op_bot_7')
// (4, 11, 'sp4_v_b_3')
// (5, 7, 'sp4_h_r_14')
// (5, 9, 'neigh_op_tnl_7')
// (5, 10, 'neigh_op_lft_7')
// (5, 11, 'neigh_op_bnl_7')
// (6, 7, 'local_g2_3')
// (6, 7, 'local_g3_3')
// (6, 7, 'lutff_0/in_3')
// (6, 7, 'lutff_3/in_3')
// (6, 7, 'sp4_h_r_27')
// (7, 7, 'sp4_h_r_38')
// (8, 7, 'sp4_h_l_38')

wire n134;
// (3, 9, 'neigh_op_tnr_3')
// (3, 10, 'neigh_op_rgt_3')
// (3, 11, 'neigh_op_bnr_3')
// (4, 9, 'neigh_op_top_3')
// (4, 10, 'local_g1_3')
// (4, 10, 'lutff_3/out')
// (4, 10, 'lutff_7/in_1')
// (4, 11, 'local_g1_3')
// (4, 11, 'lutff_3/in_1')
// (4, 11, 'neigh_op_bot_3')
// (5, 9, 'neigh_op_tnl_3')
// (5, 10, 'neigh_op_lft_3')
// (5, 11, 'neigh_op_bnl_3')

wire n135;
// (3, 9, 'sp12_h_r_1')
// (4, 9, 'sp12_h_r_2')
// (5, 9, 'sp12_h_r_5')
// (6, 9, 'sp12_h_r_6')
// (7, 8, 'neigh_op_tnr_1')
// (7, 9, 'neigh_op_rgt_1')
// (7, 9, 'sp12_h_r_9')
// (7, 10, 'neigh_op_bnr_1')
// (8, 8, 'neigh_op_top_1')
// (8, 9, 'local_g1_2')
// (8, 9, 'lutff_0/in_3')
// (8, 9, 'lutff_1/out')
// (8, 9, 'sp12_h_r_10')
// (8, 10, 'neigh_op_bot_1')
// (9, 8, 'neigh_op_tnl_1')
// (9, 9, 'neigh_op_lft_1')
// (9, 9, 'sp12_h_r_13')
// (9, 10, 'neigh_op_bnl_1')
// (10, 9, 'sp12_h_r_14')
// (11, 9, 'sp12_h_r_17')
// (12, 9, 'sp12_h_r_18')
// (13, 9, 'span12_horz_18')

wire n136;
// (3, 9, 'sp4_h_r_8')
// (4, 8, 'neigh_op_tnr_0')
// (4, 9, 'neigh_op_rgt_0')
// (4, 9, 'sp4_h_r_21')
// (4, 10, 'neigh_op_bnr_0')
// (5, 6, 'sp4_r_v_b_36')
// (5, 7, 'sp4_r_v_b_25')
// (5, 8, 'neigh_op_top_0')
// (5, 8, 'sp4_r_v_b_12')
// (5, 9, 'lutff_0/out')
// (5, 9, 'sp4_h_r_32')
// (5, 9, 'sp4_r_v_b_1')
// (5, 10, 'neigh_op_bot_0')
// (6, 5, 'sp4_v_t_36')
// (6, 6, 'local_g2_4')
// (6, 6, 'lutff_5/in_3')
// (6, 6, 'lutff_7/in_3')
// (6, 6, 'sp4_r_v_b_45')
// (6, 6, 'sp4_v_b_36')
// (6, 7, 'local_g0_3')
// (6, 7, 'lutff_3/in_2')
// (6, 7, 'sp4_r_v_b_32')
// (6, 7, 'sp4_v_b_25')
// (6, 8, 'neigh_op_tnl_0')
// (6, 8, 'sp4_r_v_b_21')
// (6, 8, 'sp4_v_b_12')
// (6, 9, 'neigh_op_lft_0')
// (6, 9, 'sp4_h_r_45')
// (6, 9, 'sp4_r_v_b_8')
// (6, 9, 'sp4_v_b_1')
// (6, 10, 'neigh_op_bnl_0')
// (7, 5, 'sp4_v_t_45')
// (7, 6, 'local_g2_5')
// (7, 6, 'lutff_3/in_2')
// (7, 6, 'sp4_v_b_45')
// (7, 7, 'sp4_v_b_32')
// (7, 8, 'sp4_v_b_21')
// (7, 9, 'sp4_h_l_45')
// (7, 9, 'sp4_v_b_8')

wire n137;
// (3, 10, 'neigh_op_tnr_0')
// (3, 11, 'neigh_op_rgt_0')
// (3, 12, 'neigh_op_bnr_0')
// (4, 8, 'sp4_r_v_b_36')
// (4, 9, 'sp4_r_v_b_25')
// (4, 10, 'neigh_op_top_0')
// (4, 10, 'sp4_r_v_b_12')
// (4, 11, 'local_g1_1')
// (4, 11, 'lutff_0/out')
// (4, 11, 'lutff_1/in_3')
// (4, 11, 'sp4_r_v_b_1')
// (4, 12, 'neigh_op_bot_0')
// (5, 7, 'sp4_v_t_36')
// (5, 8, 'sp4_v_b_36')
// (5, 9, 'sp4_v_b_25')
// (5, 10, 'neigh_op_tnl_0')
// (5, 10, 'sp4_v_b_12')
// (5, 11, 'neigh_op_lft_0')
// (5, 11, 'sp4_v_b_1')
// (5, 12, 'neigh_op_bnl_0')

wire n138;
// (3, 10, 'neigh_op_tnr_1')
// (3, 11, 'neigh_op_rgt_1')
// (3, 12, 'neigh_op_bnr_1')
// (4, 10, 'local_g1_1')
// (4, 10, 'lutff_7/in_3')
// (4, 10, 'neigh_op_top_1')
// (4, 11, 'lutff_1/out')
// (4, 12, 'neigh_op_bot_1')
// (5, 10, 'neigh_op_tnl_1')
// (5, 11, 'neigh_op_lft_1')
// (5, 12, 'neigh_op_bnl_1')

reg n139 = 0;
// (3, 10, 'neigh_op_tnr_3')
// (3, 11, 'neigh_op_rgt_3')
// (3, 12, 'neigh_op_bnr_3')
// (4, 10, 'neigh_op_top_3')
// (4, 11, 'local_g0_3')
// (4, 11, 'lutff_3/out')
// (4, 11, 'lutff_7/in_0')
// (4, 12, 'neigh_op_bot_3')
// (5, 10, 'neigh_op_tnl_3')
// (5, 11, 'neigh_op_lft_3')
// (5, 12, 'neigh_op_bnl_3')

reg n140 = 0;
// (3, 10, 'neigh_op_tnr_4')
// (3, 11, 'neigh_op_rgt_4')
// (3, 12, 'neigh_op_bnr_4')
// (4, 10, 'neigh_op_top_4')
// (4, 11, 'local_g0_4')
// (4, 11, 'lutff_4/out')
// (4, 11, 'lutff_6/in_0')
// (4, 12, 'neigh_op_bot_4')
// (5, 10, 'neigh_op_tnl_4')
// (5, 11, 'neigh_op_lft_4')
// (5, 12, 'neigh_op_bnl_4')

reg n141 = 0;
// (3, 10, 'neigh_op_tnr_7')
// (3, 11, 'neigh_op_rgt_7')
// (3, 12, 'neigh_op_bnr_7')
// (4, 10, 'neigh_op_top_7')
// (4, 11, 'local_g1_7')
// (4, 11, 'lutff_4/in_0')
// (4, 11, 'lutff_7/out')
// (4, 12, 'neigh_op_bot_7')
// (5, 10, 'neigh_op_tnl_7')
// (5, 11, 'neigh_op_lft_7')
// (5, 12, 'neigh_op_bnl_7')

reg n142 = 0;
// (3, 11, 'neigh_op_tnr_2')
// (3, 12, 'neigh_op_rgt_2')
// (3, 13, 'neigh_op_bnr_2')
// (4, 11, 'local_g0_2')
// (4, 11, 'lutff_0/in_0')
// (4, 11, 'neigh_op_top_2')
// (4, 12, 'local_g1_2')
// (4, 12, 'lutff_2/out')
// (4, 12, 'lutff_6/in_1')
// (4, 13, 'neigh_op_bot_2')
// (5, 11, 'neigh_op_tnl_2')
// (5, 12, 'neigh_op_lft_2')
// (5, 13, 'neigh_op_bnl_2')

reg n143 = 0;
// (3, 11, 'neigh_op_tnr_3')
// (3, 12, 'neigh_op_rgt_3')
// (3, 13, 'neigh_op_bnr_3')
// (4, 11, 'neigh_op_top_3')
// (4, 12, 'local_g0_3')
// (4, 12, 'lutff_3/out')
// (4, 12, 'lutff_7/in_0')
// (4, 13, 'neigh_op_bot_3')
// (5, 11, 'neigh_op_tnl_3')
// (5, 12, 'neigh_op_lft_3')
// (5, 13, 'neigh_op_bnl_3')

reg n144 = 0;
// (3, 11, 'neigh_op_tnr_6')
// (3, 12, 'neigh_op_rgt_6')
// (3, 13, 'neigh_op_bnr_6')
// (4, 11, 'neigh_op_top_6')
// (4, 12, 'local_g1_6')
// (4, 12, 'lutff_3/in_0')
// (4, 12, 'lutff_6/out')
// (4, 13, 'neigh_op_bot_6')
// (5, 11, 'neigh_op_tnl_6')
// (5, 12, 'neigh_op_lft_6')
// (5, 13, 'neigh_op_bnl_6')

reg n145 = 0;
// (3, 11, 'neigh_op_tnr_7')
// (3, 12, 'neigh_op_rgt_7')
// (3, 13, 'neigh_op_bnr_7')
// (4, 11, 'neigh_op_top_7')
// (4, 12, 'local_g2_7')
// (4, 12, 'lutff_1/in_0')
// (4, 12, 'lutff_7/out')
// (4, 13, 'neigh_op_bot_7')
// (5, 11, 'neigh_op_tnl_7')
// (5, 12, 'neigh_op_lft_7')
// (5, 13, 'neigh_op_bnl_7')

reg n146 = 0;
// (3, 12, 'neigh_op_tnr_5')
// (3, 13, 'neigh_op_rgt_5')
// (3, 14, 'neigh_op_bnr_5')
// (4, 12, 'neigh_op_top_5')
// (4, 13, 'local_g1_5')
// (4, 13, 'lutff_5/out')
// (4, 13, 'lutff_6/in_0')
// (4, 14, 'neigh_op_bot_5')
// (5, 12, 'neigh_op_tnl_5')
// (5, 13, 'neigh_op_lft_5')
// (5, 14, 'neigh_op_bnl_5')

reg n147 = 0;
// (3, 12, 'neigh_op_tnr_6')
// (3, 13, 'neigh_op_rgt_6')
// (3, 14, 'neigh_op_bnr_6')
// (4, 12, 'neigh_op_top_6')
// (4, 13, 'local_g1_6')
// (4, 13, 'lutff_1/in_0')
// (4, 13, 'lutff_6/out')
// (4, 14, 'neigh_op_bot_6')
// (5, 12, 'neigh_op_tnl_6')
// (5, 13, 'neigh_op_lft_6')
// (5, 14, 'neigh_op_bnl_6')

reg n148 = 0;
// (3, 12, 'sp12_h_r_0')
// (4, 12, 'sp12_h_r_3')
// (5, 12, 'sp12_h_r_4')
// (6, 12, 'sp12_h_r_7')
// (7, 12, 'sp12_h_r_8')
// (8, 11, 'neigh_op_tnr_2')
// (8, 12, 'neigh_op_rgt_2')
// (8, 12, 'sp12_h_r_11')
// (8, 13, 'neigh_op_bnr_2')
// (9, 11, 'neigh_op_top_2')
// (9, 12, 'lutff_2/out')
// (9, 12, 'sp12_h_r_12')
// (9, 13, 'neigh_op_bot_2')
// (10, 11, 'neigh_op_tnl_2')
// (10, 12, 'neigh_op_lft_2')
// (10, 12, 'sp12_h_r_15')
// (10, 13, 'neigh_op_bnl_2')
// (11, 12, 'local_g0_0')
// (11, 12, 'lutff_2/in_0')
// (11, 12, 'sp12_h_r_16')
// (12, 12, 'sp12_h_r_19')
// (13, 12, 'span12_horz_19')

wire n149;
// (3, 12, 'sp4_h_r_0')
// (4, 7, 'sp4_r_v_b_43')
// (4, 8, 'sp4_r_v_b_30')
// (4, 9, 'sp4_r_v_b_19')
// (4, 10, 'sp4_r_v_b_6')
// (4, 11, 'neigh_op_tnr_4')
// (4, 12, 'neigh_op_rgt_4')
// (4, 12, 'sp4_h_r_13')
// (4, 13, 'neigh_op_bnr_4')
// (5, 4, 'sp12_v_t_23')
// (5, 5, 'local_g2_7')
// (5, 5, 'lutff_2/in_3')
// (5, 5, 'lutff_4/in_1')
// (5, 5, 'sp12_v_b_23')
// (5, 5, 'sp4_r_v_b_37')
// (5, 6, 'sp12_v_b_20')
// (5, 6, 'sp4_h_r_11')
// (5, 6, 'sp4_r_v_b_24')
// (5, 6, 'sp4_v_t_43')
// (5, 7, 'sp12_v_b_19')
// (5, 7, 'sp4_r_v_b_13')
// (5, 7, 'sp4_v_b_43')
// (5, 8, 'sp12_v_b_16')
// (5, 8, 'sp4_r_v_b_0')
// (5, 8, 'sp4_v_b_30')
// (5, 9, 'sp12_v_b_15')
// (5, 9, 'sp4_r_v_b_44')
// (5, 9, 'sp4_v_b_19')
// (5, 10, 'sp12_v_b_12')
// (5, 10, 'sp4_r_v_b_33')
// (5, 10, 'sp4_v_b_6')
// (5, 11, 'neigh_op_top_4')
// (5, 11, 'sp12_v_b_11')
// (5, 11, 'sp4_r_v_b_20')
// (5, 12, 'lutff_4/out')
// (5, 12, 'sp12_v_b_8')
// (5, 12, 'sp4_h_r_24')
// (5, 12, 'sp4_r_v_b_9')
// (5, 13, 'neigh_op_bot_4')
// (5, 13, 'sp12_v_b_7')
// (5, 14, 'sp12_v_b_4')
// (5, 15, 'sp12_v_b_3')
// (5, 16, 'sp12_v_b_0')
// (6, 4, 'sp4_v_t_37')
// (6, 5, 'sp4_r_v_b_44')
// (6, 5, 'sp4_v_b_37')
// (6, 6, 'local_g0_6')
// (6, 6, 'local_g1_6')
// (6, 6, 'lutff_1/in_3')
// (6, 6, 'lutff_4/in_3')
// (6, 6, 'lutff_5/in_2')
// (6, 6, 'lutff_7/in_2')
// (6, 6, 'sp4_h_r_22')
// (6, 6, 'sp4_r_v_b_33')
// (6, 6, 'sp4_v_b_24')
// (6, 7, 'local_g1_5')
// (6, 7, 'lutff_3/in_1')
// (6, 7, 'sp4_r_v_b_20')
// (6, 7, 'sp4_v_b_13')
// (6, 8, 'sp4_r_v_b_9')
// (6, 8, 'sp4_v_b_0')
// (6, 8, 'sp4_v_t_44')
// (6, 9, 'sp4_r_v_b_43')
// (6, 9, 'sp4_v_b_44')
// (6, 10, 'sp4_r_v_b_30')
// (6, 10, 'sp4_v_b_33')
// (6, 11, 'neigh_op_tnl_4')
// (6, 11, 'sp4_r_v_b_19')
// (6, 11, 'sp4_v_b_20')
// (6, 12, 'neigh_op_lft_4')
// (6, 12, 'sp4_h_r_37')
// (6, 12, 'sp4_r_v_b_6')
// (6, 12, 'sp4_v_b_9')
// (6, 13, 'neigh_op_bnl_4')
// (7, 4, 'sp4_v_t_44')
// (7, 5, 'local_g2_4')
// (7, 5, 'lutff_4/in_2')
// (7, 5, 'sp4_v_b_44')
// (7, 6, 'local_g3_3')
// (7, 6, 'lutff_0/in_2')
// (7, 6, 'lutff_2/in_2')
// (7, 6, 'lutff_6/in_2')
// (7, 6, 'sp4_h_r_35')
// (7, 6, 'sp4_v_b_33')
// (7, 7, 'sp4_v_b_20')
// (7, 8, 'sp4_v_b_9')
// (7, 8, 'sp4_v_t_43')
// (7, 9, 'sp4_v_b_43')
// (7, 10, 'sp4_v_b_30')
// (7, 11, 'sp4_v_b_19')
// (7, 12, 'sp4_h_l_37')
// (7, 12, 'sp4_v_b_6')
// (8, 6, 'sp4_h_r_46')
// (9, 6, 'sp4_h_l_46')

reg n150 = 0;
// (3, 13, 'neigh_op_tnr_6')
// (3, 14, 'neigh_op_rgt_6')
// (3, 15, 'neigh_op_bnr_6')
// (4, 13, 'neigh_op_top_6')
// (4, 14, 'local_g1_6')
// (4, 14, 'lutff_1/in_0')
// (4, 14, 'lutff_6/out')
// (4, 15, 'neigh_op_bot_6')
// (5, 13, 'neigh_op_tnl_6')
// (5, 14, 'neigh_op_lft_6')
// (5, 15, 'neigh_op_bnl_6')

wire n151;
// (4, 1, 'neigh_op_tnr_1')
// (4, 2, 'neigh_op_rgt_1')
// (4, 3, 'neigh_op_bnr_1')
// (5, 1, 'neigh_op_top_1')
// (5, 2, 'local_g1_1')
// (5, 2, 'local_g2_1')
// (5, 2, 'lutff_1/out')
// (5, 2, 'lutff_4/in_3')
// (5, 2, 'lutff_6/in_2')
// (5, 3, 'neigh_op_bot_1')
// (6, 1, 'neigh_op_tnl_1')
// (6, 2, 'neigh_op_lft_1')
// (6, 3, 'neigh_op_bnl_1')

wire n152;
// (4, 1, 'neigh_op_tnr_2')
// (4, 2, 'neigh_op_rgt_2')
// (4, 3, 'neigh_op_bnr_2')
// (5, 1, 'neigh_op_top_2')
// (5, 2, 'local_g0_2')
// (5, 2, 'lutff_2/out')
// (5, 2, 'lutff_5/in_3')
// (5, 3, 'neigh_op_bot_2')
// (6, 1, 'neigh_op_tnl_2')
// (6, 2, 'neigh_op_lft_2')
// (6, 3, 'neigh_op_bnl_2')

wire n153;
// (4, 1, 'neigh_op_tnr_4')
// (4, 2, 'neigh_op_rgt_4')
// (4, 3, 'neigh_op_bnr_4')
// (5, 1, 'neigh_op_top_4')
// (5, 2, 'local_g2_4')
// (5, 2, 'lutff_4/out')
// (5, 2, 'lutff_7/in_1')
// (5, 3, 'neigh_op_bot_4')
// (6, 1, 'neigh_op_tnl_4')
// (6, 2, 'neigh_op_lft_4')
// (6, 3, 'neigh_op_bnl_4')

wire n154;
// (4, 1, 'neigh_op_tnr_6')
// (4, 2, 'neigh_op_rgt_6')
// (4, 3, 'neigh_op_bnr_6')
// (5, 1, 'neigh_op_top_6')
// (5, 2, 'lutff_6/out')
// (5, 3, 'neigh_op_bot_6')
// (6, 1, 'neigh_op_tnl_6')
// (6, 2, 'neigh_op_lft_6')
// (6, 3, 'local_g2_6')
// (6, 3, 'lutff_0/in_2')
// (6, 3, 'neigh_op_bnl_6')

wire n155;
// (4, 1, 'neigh_op_tnr_7')
// (4, 2, 'neigh_op_rgt_7')
// (4, 3, 'neigh_op_bnr_7')
// (5, 1, 'neigh_op_top_7')
// (5, 1, 'sp4_r_v_b_26')
// (5, 2, 'lutff_7/out')
// (5, 2, 'sp4_r_v_b_15')
// (5, 3, 'neigh_op_bot_7')
// (5, 3, 'sp4_r_v_b_2')
// (6, 0, 'span4_vert_26')
// (6, 1, 'neigh_op_tnl_7')
// (6, 1, 'sp4_v_b_26')
// (6, 2, 'neigh_op_lft_7')
// (6, 2, 'sp4_v_b_15')
// (6, 3, 'neigh_op_bnl_7')
// (6, 3, 'sp4_h_r_8')
// (6, 3, 'sp4_v_b_2')
// (7, 3, 'local_g1_5')
// (7, 3, 'lutff_7/in_1')
// (7, 3, 'sp4_h_r_21')
// (8, 3, 'sp4_h_r_32')
// (9, 3, 'sp4_h_r_45')
// (10, 3, 'sp4_h_l_45')

wire n156;
// (4, 2, 'neigh_op_tnr_1')
// (4, 3, 'neigh_op_rgt_1')
// (4, 4, 'neigh_op_bnr_1')
// (5, 2, 'neigh_op_top_1')
// (5, 3, 'lutff_1/out')
// (5, 4, 'neigh_op_bot_1')
// (6, 2, 'neigh_op_tnl_1')
// (6, 3, 'neigh_op_lft_1')
// (6, 4, 'local_g3_1')
// (6, 4, 'lutff_4/in_2')
// (6, 4, 'neigh_op_bnl_1')

wire n157;
// (4, 2, 'neigh_op_tnr_2')
// (4, 3, 'neigh_op_rgt_2')
// (4, 4, 'neigh_op_bnr_2')
// (5, 1, 'sp4_r_v_b_45')
// (5, 2, 'neigh_op_top_2')
// (5, 2, 'sp4_r_v_b_32')
// (5, 3, 'local_g1_2')
// (5, 3, 'lutff_2/out')
// (5, 3, 'lutff_7/in_2')
// (5, 3, 'sp4_r_v_b_21')
// (5, 4, 'local_g0_2')
// (5, 4, 'lutff_6/in_2')
// (5, 4, 'neigh_op_bot_2')
// (5, 4, 'sp4_r_v_b_8')
// (6, 0, 'span4_vert_45')
// (6, 1, 'sp4_v_b_45')
// (6, 2, 'neigh_op_tnl_2')
// (6, 2, 'sp4_v_b_32')
// (6, 3, 'neigh_op_lft_2')
// (6, 3, 'sp4_v_b_21')
// (6, 4, 'neigh_op_bnl_2')
// (6, 4, 'sp4_h_r_8')
// (6, 4, 'sp4_v_b_8')
// (7, 4, 'local_g0_5')
// (7, 4, 'lutff_1/in_0')
// (7, 4, 'sp4_h_r_21')
// (8, 4, 'sp4_h_r_32')
// (9, 4, 'sp4_h_r_45')
// (10, 4, 'sp4_h_l_45')

wire n158;
// (4, 2, 'neigh_op_tnr_3')
// (4, 3, 'neigh_op_rgt_3')
// (4, 4, 'neigh_op_bnr_3')
// (5, 2, 'neigh_op_top_3')
// (5, 3, 'local_g1_3')
// (5, 3, 'lutff_3/out')
// (5, 3, 'lutff_6/in_2')
// (5, 4, 'neigh_op_bot_3')
// (6, 2, 'neigh_op_tnl_3')
// (6, 3, 'neigh_op_lft_3')
// (6, 4, 'neigh_op_bnl_3')

wire n159;
// (4, 2, 'neigh_op_tnr_5')
// (4, 3, 'neigh_op_rgt_5')
// (4, 4, 'neigh_op_bnr_5')
// (5, 2, 'neigh_op_top_5')
// (5, 3, 'local_g1_5')
// (5, 3, 'lutff_3/in_3')
// (5, 3, 'lutff_5/out')
// (5, 4, 'neigh_op_bot_5')
// (6, 2, 'neigh_op_tnl_5')
// (6, 3, 'neigh_op_lft_5')
// (6, 4, 'neigh_op_bnl_5')

wire n160;
// (4, 2, 'neigh_op_tnr_6')
// (4, 2, 'sp4_r_v_b_41')
// (4, 3, 'neigh_op_rgt_6')
// (4, 3, 'sp4_r_v_b_28')
// (4, 4, 'neigh_op_bnr_6')
// (4, 4, 'sp4_r_v_b_17')
// (4, 5, 'sp4_r_v_b_4')
// (4, 6, 'sp4_r_v_b_37')
// (4, 7, 'sp4_r_v_b_24')
// (4, 8, 'sp4_r_v_b_13')
// (4, 9, 'sp4_r_v_b_0')
// (5, 1, 'sp4_v_t_41')
// (5, 2, 'neigh_op_top_6')
// (5, 2, 'sp4_v_b_41')
// (5, 3, 'lutff_6/out')
// (5, 3, 'sp4_v_b_28')
// (5, 4, 'neigh_op_bot_6')
// (5, 4, 'sp4_v_b_17')
// (5, 5, 'sp4_v_b_4')
// (5, 5, 'sp4_v_t_37')
// (5, 6, 'sp4_v_b_37')
// (5, 7, 'sp4_v_b_24')
// (5, 8, 'sp4_v_b_13')
// (5, 9, 'local_g0_0')
// (5, 9, 'lutff_2/in_2')
// (5, 9, 'sp4_v_b_0')
// (6, 2, 'neigh_op_tnl_6')
// (6, 3, 'neigh_op_lft_6')
// (6, 4, 'neigh_op_bnl_6')

reg \d_out[5] = 0 ;
// (4, 2, 'neigh_op_tnr_7')
// (4, 3, 'neigh_op_rgt_7')
// (4, 4, 'neigh_op_bnr_7')
// (5, 0, 'io_0/D_OUT_0')
// (5, 0, 'io_0/PAD')
// (5, 0, 'local_g0_2')
// (5, 0, 'span12_vert_18')
// (5, 1, 'sp12_v_b_18')
// (5, 2, 'neigh_op_top_7')
// (5, 2, 'sp12_v_b_17')
// (5, 3, 'lutff_7/out')
// (5, 3, 'sp12_v_b_14')
// (5, 4, 'neigh_op_bot_7')
// (5, 4, 'sp12_v_b_13')
// (5, 5, 'sp12_v_b_10')
// (5, 6, 'sp12_v_b_9')
// (5, 7, 'sp12_v_b_6')
// (5, 8, 'sp12_v_b_5')
// (5, 9, 'sp12_v_b_2')
// (5, 10, 'sp12_v_b_1')
// (6, 2, 'neigh_op_tnl_7')
// (6, 3, 'neigh_op_lft_7')
// (6, 4, 'neigh_op_bnl_7')

wire n162;
// (4, 2, 'sp4_h_r_9')
// (5, 2, 'sp4_h_r_20')
// (6, 2, 'local_g2_1')
// (6, 2, 'lutff_5/in_2')
// (6, 2, 'sp4_h_r_33')
// (7, 1, 'local_g1_6')
// (7, 1, 'lutff_0/in_3')
// (7, 1, 'lutff_1/in_2')
// (7, 1, 'sp4_r_v_b_30')
// (7, 2, 'local_g2_3')
// (7, 2, 'lutff_2/in_3')
// (7, 2, 'neigh_op_tnr_3')
// (7, 2, 'sp4_h_r_44')
// (7, 2, 'sp4_r_v_b_19')
// (7, 3, 'neigh_op_rgt_3')
// (7, 3, 'sp4_r_v_b_38')
// (7, 3, 'sp4_r_v_b_6')
// (7, 4, 'neigh_op_bnr_3')
// (7, 4, 'sp4_r_v_b_27')
// (7, 5, 'sp4_r_v_b_14')
// (7, 6, 'sp4_r_v_b_3')
// (8, 0, 'span4_vert_30')
// (8, 1, 'sp4_v_b_30')
// (8, 2, 'local_g1_3')
// (8, 2, 'lutff_0/in_2')
// (8, 2, 'neigh_op_top_3')
// (8, 2, 'sp4_h_l_44')
// (8, 2, 'sp4_v_b_19')
// (8, 2, 'sp4_v_t_38')
// (8, 3, 'lutff_3/out')
// (8, 3, 'sp4_v_b_38')
// (8, 3, 'sp4_v_b_6')
// (8, 4, 'neigh_op_bot_3')
// (8, 4, 'sp4_v_b_27')
// (8, 5, 'sp4_v_b_14')
// (8, 6, 'sp4_v_b_3')
// (9, 2, 'neigh_op_tnl_3')
// (9, 3, 'neigh_op_lft_3')
// (9, 4, 'neigh_op_bnl_3')

reg n163 = 0;
// (4, 3, 'neigh_op_tnr_2')
// (4, 4, 'neigh_op_rgt_2')
// (4, 5, 'neigh_op_bnr_2')
// (5, 2, 'sp4_r_v_b_45')
// (5, 3, 'local_g0_3')
// (5, 3, 'lutff_2/in_3')
// (5, 3, 'neigh_op_top_2')
// (5, 3, 'sp4_r_v_b_32')
// (5, 4, 'lutff_2/out')
// (5, 4, 'sp4_r_v_b_21')
// (5, 5, 'neigh_op_bot_2')
// (5, 5, 'sp4_r_v_b_8')
// (6, 1, 'sp4_v_t_45')
// (6, 2, 'sp4_v_b_45')
// (6, 3, 'neigh_op_tnl_2')
// (6, 3, 'sp4_v_b_32')
// (6, 4, 'neigh_op_lft_2')
// (6, 4, 'sp4_v_b_21')
// (6, 5, 'neigh_op_bnl_2')
// (6, 5, 'sp4_v_b_8')

reg n164 = 0;
// (4, 3, 'neigh_op_tnr_4')
// (4, 4, 'neigh_op_rgt_4')
// (4, 5, 'neigh_op_bnr_4')
// (5, 3, 'neigh_op_top_4')
// (5, 4, 'local_g1_4')
// (5, 4, 'lutff_4/out')
// (5, 4, 'lutff_7/in_0')
// (5, 5, 'neigh_op_bot_4')
// (6, 3, 'neigh_op_tnl_4')
// (6, 4, 'neigh_op_lft_4')
// (6, 5, 'neigh_op_bnl_4')

reg n165 = 0;
// (4, 3, 'neigh_op_tnr_6')
// (4, 4, 'neigh_op_rgt_6')
// (4, 5, 'neigh_op_bnr_6')
// (5, 3, 'neigh_op_top_6')
// (5, 4, 'local_g0_6')
// (5, 4, 'lutff_4/in_0')
// (5, 4, 'lutff_6/out')
// (5, 5, 'neigh_op_bot_6')
// (6, 3, 'neigh_op_tnl_6')
// (6, 4, 'neigh_op_lft_6')
// (6, 5, 'neigh_op_bnl_6')

reg n166 = 0;
// (4, 3, 'neigh_op_tnr_7')
// (4, 4, 'neigh_op_rgt_7')
// (4, 5, 'neigh_op_bnr_7')
// (5, 3, 'neigh_op_top_7')
// (5, 4, 'local_g1_7')
// (5, 4, 'lutff_2/in_0')
// (5, 4, 'lutff_7/out')
// (5, 5, 'neigh_op_bot_7')
// (6, 3, 'neigh_op_tnl_7')
// (6, 4, 'neigh_op_lft_7')
// (6, 5, 'neigh_op_bnl_7')

wire n167;
// (4, 3, 'sp4_h_r_0')
// (5, 3, 'local_g0_5')
// (5, 3, 'lutff_6/in_1')
// (5, 3, 'sp4_h_r_13')
// (6, 1, 'neigh_op_tnr_6')
// (6, 2, 'neigh_op_rgt_6')
// (6, 3, 'local_g1_6')
// (6, 3, 'lutff_2/in_1')
// (6, 3, 'neigh_op_bnr_6')
// (6, 3, 'sp4_h_r_24')
// (7, 1, 'neigh_op_top_6')
// (7, 1, 'sp4_r_v_b_24')
// (7, 2, 'lutff_6/out')
// (7, 2, 'sp4_r_v_b_13')
// (7, 3, 'local_g1_6')
// (7, 3, 'lutff_7/in_2')
// (7, 3, 'neigh_op_bot_6')
// (7, 3, 'sp4_h_r_37')
// (7, 3, 'sp4_r_v_b_0')
// (8, 0, 'span4_vert_24')
// (8, 1, 'neigh_op_tnl_6')
// (8, 1, 'sp4_v_b_24')
// (8, 2, 'neigh_op_lft_6')
// (8, 2, 'sp4_v_b_13')
// (8, 3, 'neigh_op_bnl_6')
// (8, 3, 'sp4_h_l_37')
// (8, 3, 'sp4_v_b_0')

wire n168;
// (4, 3, 'sp4_r_v_b_42')
// (4, 4, 'neigh_op_tnr_1')
// (4, 4, 'sp4_r_v_b_31')
// (4, 5, 'neigh_op_rgt_1')
// (4, 5, 'sp4_r_v_b_18')
// (4, 6, 'neigh_op_bnr_1')
// (4, 6, 'sp4_r_v_b_7')
// (5, 2, 'sp4_v_t_42')
// (5, 3, 'sp4_v_b_42')
// (5, 4, 'neigh_op_top_1')
// (5, 4, 'sp4_v_b_31')
// (5, 5, 'local_g0_1')
// (5, 5, 'lutff_1/out')
// (5, 5, 'lutff_5/in_2')
// (5, 5, 'sp4_v_b_18')
// (5, 6, 'local_g0_7')
// (5, 6, 'lutff_0/in_3')
// (5, 6, 'neigh_op_bot_1')
// (5, 6, 'sp4_v_b_7')
// (6, 4, 'neigh_op_tnl_1')
// (6, 5, 'neigh_op_lft_1')
// (6, 6, 'neigh_op_bnl_1')

wire n169;
// (4, 3, 'sp4_r_v_b_45')
// (4, 4, 'sp4_r_v_b_32')
// (4, 5, 'sp4_r_v_b_21')
// (4, 6, 'sp4_r_v_b_8')
// (5, 2, 'sp4_v_t_45')
// (5, 3, 'sp4_v_b_45')
// (5, 4, 'sp4_v_b_32')
// (5, 5, 'local_g1_5')
// (5, 5, 'lutff_1/in_1')
// (5, 5, 'lutff_3/in_1')
// (5, 5, 'lutff_6/in_2')
// (5, 5, 'sp4_v_b_21')
// (5, 6, 'sp4_h_r_8')
// (5, 6, 'sp4_v_b_8')
// (6, 5, 'neigh_op_tnr_0')
// (6, 6, 'local_g2_0')
// (6, 6, 'local_g3_0')
// (6, 6, 'lutff_0/in_3')
// (6, 6, 'lutff_3/in_2')
// (6, 6, 'lutff_6/in_2')
// (6, 6, 'neigh_op_rgt_0')
// (6, 6, 'sp4_h_r_21')
// (6, 7, 'neigh_op_bnr_0')
// (7, 5, 'local_g1_0')
// (7, 5, 'lutff_4/in_3')
// (7, 5, 'neigh_op_top_0')
// (7, 6, 'local_g1_0')
// (7, 6, 'lutff_0/out')
// (7, 6, 'lutff_6/in_1')
// (7, 6, 'sp4_h_r_32')
// (7, 7, 'neigh_op_bot_0')
// (8, 5, 'neigh_op_tnl_0')
// (8, 6, 'neigh_op_lft_0')
// (8, 6, 'sp4_h_r_45')
// (8, 7, 'neigh_op_bnl_0')
// (9, 6, 'sp4_h_l_45')

wire n170;
// (4, 4, 'neigh_op_tnr_0')
// (4, 5, 'neigh_op_rgt_0')
// (4, 6, 'neigh_op_bnr_0')
// (4, 6, 'sp4_r_v_b_41')
// (4, 7, 'sp4_r_v_b_28')
// (4, 8, 'local_g2_7')
// (4, 8, 'local_g3_1')
// (4, 8, 'lutff_5/in_3')
// (4, 8, 'lutff_6/in_3')
// (4, 8, 'lutff_7/in_3')
// (4, 8, 'sp4_r_v_b_17')
// (4, 8, 'sp4_r_v_b_39')
// (4, 9, 'sp4_r_v_b_26')
// (4, 9, 'sp4_r_v_b_4')
// (4, 10, 'sp4_r_v_b_15')
// (4, 11, 'sp4_r_v_b_2')
// (5, 1, 'sp12_v_t_23')
// (5, 2, 'sp12_v_b_23')
// (5, 2, 'sp4_r_v_b_36')
// (5, 3, 'local_g1_1')
// (5, 3, 'lutff_7/in_3')
// (5, 3, 'sp12_v_b_20')
// (5, 3, 'sp4_r_v_b_25')
// (5, 4, 'neigh_op_top_0')
// (5, 4, 'sp12_v_b_19')
// (5, 4, 'sp4_r_v_b_12')
// (5, 4, 'sp4_r_v_b_44')
// (5, 5, 'lutff_0/out')
// (5, 5, 'sp12_v_b_16')
// (5, 5, 'sp4_r_v_b_1')
// (5, 5, 'sp4_r_v_b_33')
// (5, 5, 'sp4_v_t_41')
// (5, 6, 'neigh_op_bot_0')
// (5, 6, 'sp12_v_b_15')
// (5, 6, 'sp4_r_v_b_20')
// (5, 6, 'sp4_v_b_41')
// (5, 7, 'sp12_v_b_12')
// (5, 7, 'sp4_r_v_b_9')
// (5, 7, 'sp4_v_b_28')
// (5, 7, 'sp4_v_t_39')
// (5, 8, 'local_g2_3')
// (5, 8, 'lutff_2/in_1')
// (5, 8, 'lutff_3/in_2')
// (5, 8, 'sp12_v_b_11')
// (5, 8, 'sp4_r_v_b_37')
// (5, 8, 'sp4_r_v_b_44')
// (5, 8, 'sp4_v_b_17')
// (5, 8, 'sp4_v_b_39')
// (5, 9, 'sp12_v_b_8')
// (5, 9, 'sp4_r_v_b_24')
// (5, 9, 'sp4_r_v_b_33')
// (5, 9, 'sp4_v_b_26')
// (5, 9, 'sp4_v_b_4')
// (5, 10, 'sp12_v_b_7')
// (5, 10, 'sp4_r_v_b_13')
// (5, 10, 'sp4_r_v_b_20')
// (5, 10, 'sp4_v_b_15')
// (5, 11, 'sp12_v_b_4')
// (5, 11, 'sp4_r_v_b_0')
// (5, 11, 'sp4_r_v_b_9')
// (5, 11, 'sp4_v_b_2')
// (5, 12, 'sp12_v_b_3')
// (5, 13, 'sp12_v_b_0')
// (6, 1, 'sp4_v_t_36')
// (6, 2, 'sp4_v_b_36')
// (6, 3, 'sp4_v_b_25')
// (6, 3, 'sp4_v_t_44')
// (6, 4, 'neigh_op_tnl_0')
// (6, 4, 'sp4_v_b_12')
// (6, 4, 'sp4_v_b_44')
// (6, 5, 'neigh_op_lft_0')
// (6, 5, 'sp4_v_b_1')
// (6, 5, 'sp4_v_b_33')
// (6, 6, 'neigh_op_bnl_0')
// (6, 6, 'sp4_v_b_20')
// (6, 7, 'sp4_v_b_9')
// (6, 7, 'sp4_v_t_37')
// (6, 7, 'sp4_v_t_44')
// (6, 8, 'sp4_v_b_37')
// (6, 8, 'sp4_v_b_44')
// (6, 9, 'sp4_v_b_24')
// (6, 9, 'sp4_v_b_33')
// (6, 10, 'local_g0_4')
// (6, 10, 'local_g0_5')
// (6, 10, 'lutff_1/in_2')
// (6, 10, 'lutff_7/in_3')
// (6, 10, 'sp4_v_b_13')
// (6, 10, 'sp4_v_b_20')
// (6, 11, 'sp4_v_b_0')
// (6, 11, 'sp4_v_b_9')

wire n171;
// (4, 4, 'neigh_op_tnr_2')
// (4, 5, 'neigh_op_rgt_2')
// (4, 5, 'sp4_r_v_b_36')
// (4, 6, 'neigh_op_bnr_2')
// (4, 6, 'sp4_r_v_b_25')
// (4, 7, 'sp4_r_v_b_12')
// (4, 8, 'sp4_r_v_b_1')
// (5, 4, 'neigh_op_top_2')
// (5, 4, 'sp4_v_t_36')
// (5, 5, 'local_g0_2')
// (5, 5, 'lutff_0/in_0')
// (5, 5, 'lutff_2/out')
// (5, 5, 'sp4_v_b_36')
// (5, 6, 'local_g0_2')
// (5, 6, 'lutff_6/in_2')
// (5, 6, 'neigh_op_bot_2')
// (5, 6, 'sp4_v_b_25')
// (5, 7, 'local_g0_4')
// (5, 7, 'lutff_0/in_2')
// (5, 7, 'sp4_v_b_12')
// (5, 8, 'sp4_v_b_1')
// (6, 4, 'neigh_op_tnl_2')
// (6, 5, 'neigh_op_lft_2')
// (6, 6, 'neigh_op_bnl_2')

wire n172;
// (4, 4, 'neigh_op_tnr_3')
// (4, 5, 'neigh_op_rgt_3')
// (4, 5, 'sp4_r_v_b_38')
// (4, 6, 'neigh_op_bnr_3')
// (4, 6, 'sp4_r_v_b_27')
// (4, 7, 'sp4_r_v_b_14')
// (4, 8, 'sp4_r_v_b_3')
// (5, 4, 'neigh_op_top_3')
// (5, 4, 'sp4_v_t_38')
// (5, 5, 'lutff_3/out')
// (5, 5, 'sp4_v_b_38')
// (5, 6, 'neigh_op_bot_3')
// (5, 6, 'sp4_v_b_27')
// (5, 7, 'sp4_v_b_14')
// (5, 8, 'local_g1_3')
// (5, 8, 'lutff_2/in_2')
// (5, 8, 'lutff_3/in_3')
// (5, 8, 'sp4_v_b_3')
// (6, 4, 'neigh_op_tnl_3')
// (6, 5, 'neigh_op_lft_3')
// (6, 6, 'neigh_op_bnl_3')

wire n173;
// (4, 4, 'neigh_op_tnr_4')
// (4, 5, 'neigh_op_rgt_4')
// (4, 6, 'neigh_op_bnr_4')
// (5, 4, 'neigh_op_top_4')
// (5, 5, 'local_g0_4')
// (5, 5, 'lutff_4/out')
// (5, 5, 'lutff_5/in_3')
// (5, 6, 'neigh_op_bot_4')
// (6, 4, 'neigh_op_tnl_4')
// (6, 5, 'neigh_op_lft_4')
// (6, 6, 'neigh_op_bnl_4')

wire n174;
// (4, 4, 'neigh_op_tnr_5')
// (4, 5, 'local_g2_5')
// (4, 5, 'lutff_3/in_2')
// (4, 5, 'neigh_op_rgt_5')
// (4, 5, 'sp4_r_v_b_42')
// (4, 6, 'neigh_op_bnr_5')
// (4, 6, 'sp4_r_v_b_31')
// (4, 7, 'sp4_r_v_b_18')
// (4, 8, 'sp4_r_v_b_7')
// (5, 2, 'sp4_r_v_b_46')
// (5, 3, 'sp4_r_v_b_35')
// (5, 4, 'neigh_op_top_5')
// (5, 4, 'sp4_r_v_b_22')
// (5, 4, 'sp4_v_t_42')
// (5, 5, 'lutff_5/out')
// (5, 5, 'sp4_r_v_b_11')
// (5, 5, 'sp4_v_b_42')
// (5, 6, 'neigh_op_bot_5')
// (5, 6, 'sp4_r_v_b_39')
// (5, 6, 'sp4_v_b_31')
// (5, 7, 'sp4_r_v_b_26')
// (5, 7, 'sp4_v_b_18')
// (5, 8, 'local_g0_7')
// (5, 8, 'lutff_0/in_3')
// (5, 8, 'lutff_4/in_3')
// (5, 8, 'sp4_r_v_b_15')
// (5, 8, 'sp4_v_b_7')
// (5, 9, 'sp4_r_v_b_2')
// (5, 10, 'sp4_r_v_b_40')
// (5, 11, 'sp4_r_v_b_29')
// (5, 12, 'sp4_r_v_b_16')
// (5, 13, 'sp4_r_v_b_5')
// (6, 1, 'sp4_v_t_46')
// (6, 2, 'sp4_v_b_46')
// (6, 3, 'sp4_v_b_35')
// (6, 4, 'neigh_op_tnl_5')
// (6, 4, 'sp4_v_b_22')
// (6, 5, 'neigh_op_lft_5')
// (6, 5, 'sp4_v_b_11')
// (6, 5, 'sp4_v_t_39')
// (6, 6, 'neigh_op_bnl_5')
// (6, 6, 'sp4_v_b_39')
// (6, 7, 'sp4_v_b_26')
// (6, 8, 'sp4_v_b_15')
// (6, 9, 'sp4_v_b_2')
// (6, 9, 'sp4_v_t_40')
// (6, 10, 'local_g2_0')
// (6, 10, 'local_g3_0')
// (6, 10, 'lutff_1/in_3')
// (6, 10, 'lutff_2/in_3')
// (6, 10, 'lutff_3/in_3')
// (6, 10, 'sp4_v_b_40')
// (6, 11, 'local_g3_5')
// (6, 11, 'lutff_1/in_3')
// (6, 11, 'lutff_5/in_3')
// (6, 11, 'sp4_v_b_29')
// (6, 12, 'sp4_v_b_16')
// (6, 13, 'sp4_v_b_5')

wire n175;
// (4, 4, 'neigh_op_tnr_6')
// (4, 5, 'neigh_op_rgt_6')
// (4, 6, 'neigh_op_bnr_6')
// (5, 4, 'neigh_op_top_6')
// (5, 5, 'local_g0_6')
// (5, 5, 'lutff_3/in_3')
// (5, 5, 'lutff_6/out')
// (5, 6, 'neigh_op_bot_6')
// (6, 4, 'neigh_op_tnl_6')
// (6, 5, 'neigh_op_lft_6')
// (6, 6, 'neigh_op_bnl_6')

reg n176 = 0;
// (4, 4, 'neigh_op_tnr_7')
// (4, 4, 'sp4_r_v_b_43')
// (4, 5, 'neigh_op_rgt_7')
// (4, 5, 'sp4_r_v_b_30')
// (4, 6, 'neigh_op_bnr_7')
// (4, 6, 'sp4_r_v_b_19')
// (4, 7, 'sp4_r_v_b_6')
// (5, 3, 'sp4_v_t_43')
// (5, 4, 'neigh_op_top_7')
// (5, 4, 'sp4_v_b_43')
// (5, 5, 'lutff_7/out')
// (5, 5, 'sp4_v_b_30')
// (5, 6, 'neigh_op_bot_7')
// (5, 6, 'sp4_v_b_19')
// (5, 7, 'local_g0_6')
// (5, 7, 'lutff_2/in_0')
// (5, 7, 'sp4_v_b_6')
// (6, 4, 'neigh_op_tnl_7')
// (6, 5, 'neigh_op_lft_7')
// (6, 6, 'neigh_op_bnl_7')

wire n177;
// (4, 4, 'sp12_h_r_1')
// (5, 4, 'sp12_h_r_2')
// (6, 4, 'sp12_h_r_5')
// (7, 4, 'sp12_h_r_6')
// (8, 3, 'neigh_op_tnr_1')
// (8, 4, 'local_g0_1')
// (8, 4, 'local_g1_1')
// (8, 4, 'lutff_2/in_2')
// (8, 4, 'lutff_4/in_1')
// (8, 4, 'neigh_op_rgt_1')
// (8, 4, 'sp12_h_r_9')
// (8, 5, 'neigh_op_bnr_1')
// (9, 3, 'neigh_op_top_1')
// (9, 4, 'lutff_1/out')
// (9, 4, 'sp12_h_r_10')
// (9, 5, 'neigh_op_bot_1')
// (10, 3, 'neigh_op_tnl_1')
// (10, 4, 'neigh_op_lft_1')
// (10, 4, 'sp12_h_r_13')
// (10, 5, 'neigh_op_bnl_1')
// (11, 4, 'sp12_h_r_14')
// (12, 4, 'sp12_h_r_17')
// (13, 4, 'span12_horz_17')

wire n178;
// (4, 5, 'neigh_op_tnr_0')
// (4, 6, 'local_g3_0')
// (4, 6, 'lutff_0/in_3')
// (4, 6, 'neigh_op_rgt_0')
// (4, 7, 'neigh_op_bnr_0')
// (4, 7, 'sp4_r_v_b_41')
// (4, 8, 'sp4_r_v_b_28')
// (4, 9, 'local_g2_7')
// (4, 9, 'local_g3_1')
// (4, 9, 'lutff_2/in_3')
// (4, 9, 'lutff_7/in_3')
// (4, 9, 'sp4_r_v_b_17')
// (4, 9, 'sp4_r_v_b_39')
// (4, 10, 'sp4_r_v_b_26')
// (4, 10, 'sp4_r_v_b_4')
// (4, 11, 'sp4_r_v_b_15')
// (4, 12, 'sp4_r_v_b_2')
// (5, 2, 'sp12_v_t_23')
// (5, 3, 'sp12_v_b_23')
// (5, 4, 'sp12_v_b_20')
// (5, 5, 'neigh_op_top_0')
// (5, 5, 'sp12_v_b_19')
// (5, 5, 'sp4_r_v_b_44')
// (5, 6, 'lutff_0/out')
// (5, 6, 'sp12_v_b_16')
// (5, 6, 'sp4_r_v_b_33')
// (5, 6, 'sp4_v_t_41')
// (5, 7, 'neigh_op_bot_0')
// (5, 7, 'sp12_v_b_15')
// (5, 7, 'sp4_r_v_b_20')
// (5, 7, 'sp4_v_b_41')
// (5, 8, 'local_g2_1')
// (5, 8, 'lutff_2/in_3')
// (5, 8, 'sp12_v_b_12')
// (5, 8, 'sp4_r_v_b_9')
// (5, 8, 'sp4_v_b_28')
// (5, 8, 'sp4_v_t_39')
// (5, 9, 'local_g3_3')
// (5, 9, 'lutff_1/in_3')
// (5, 9, 'sp12_v_b_11')
// (5, 9, 'sp4_r_v_b_37')
// (5, 9, 'sp4_v_b_17')
// (5, 9, 'sp4_v_b_39')
// (5, 10, 'sp12_v_b_8')
// (5, 10, 'sp4_r_v_b_24')
// (5, 10, 'sp4_v_b_26')
// (5, 10, 'sp4_v_b_4')
// (5, 11, 'local_g3_7')
// (5, 11, 'lutff_1/in_3')
// (5, 11, 'sp12_v_b_7')
// (5, 11, 'sp4_r_v_b_13')
// (5, 11, 'sp4_v_b_15')
// (5, 12, 'sp12_v_b_4')
// (5, 12, 'sp4_r_v_b_0')
// (5, 12, 'sp4_v_b_2')
// (5, 13, 'sp12_v_b_3')
// (5, 14, 'sp12_v_b_0')
// (6, 4, 'sp4_v_t_44')
// (6, 5, 'neigh_op_tnl_0')
// (6, 5, 'sp4_v_b_44')
// (6, 6, 'neigh_op_lft_0')
// (6, 6, 'sp4_v_b_33')
// (6, 7, 'neigh_op_bnl_0')
// (6, 7, 'sp4_v_b_20')
// (6, 8, 'sp4_v_b_9')
// (6, 8, 'sp4_v_t_37')
// (6, 9, 'sp4_v_b_37')
// (6, 10, 'sp4_v_b_24')
// (6, 11, 'local_g0_5')
// (6, 11, 'lutff_2/in_3')
// (6, 11, 'lutff_4/in_3')
// (6, 11, 'lutff_5/in_2')
// (6, 11, 'sp4_v_b_13')
// (6, 12, 'sp4_v_b_0')

wire n179;
// (4, 5, 'neigh_op_tnr_1')
// (4, 6, 'neigh_op_rgt_1')
// (4, 7, 'neigh_op_bnr_1')
// (5, 5, 'neigh_op_top_1')
// (5, 6, 'local_g2_1')
// (5, 6, 'lutff_1/out')
// (5, 6, 'lutff_3/in_2')
// (5, 6, 'lutff_6/in_1')
// (5, 7, 'neigh_op_bot_1')
// (6, 5, 'neigh_op_tnl_1')
// (6, 6, 'neigh_op_lft_1')
// (6, 7, 'neigh_op_bnl_1')

wire n180;
// (4, 5, 'neigh_op_tnr_2')
// (4, 6, 'neigh_op_rgt_2')
// (4, 7, 'neigh_op_bnr_2')
// (5, 5, 'neigh_op_top_2')
// (5, 6, 'local_g2_2')
// (5, 6, 'lutff_0/in_2')
// (5, 6, 'lutff_2/out')
// (5, 6, 'lutff_5/in_3')
// (5, 7, 'neigh_op_bot_2')
// (6, 5, 'neigh_op_tnl_2')
// (6, 6, 'neigh_op_lft_2')
// (6, 7, 'neigh_op_bnl_2')

wire n181;
// (4, 5, 'neigh_op_tnr_3')
// (4, 6, 'neigh_op_rgt_3')
// (4, 7, 'neigh_op_bnr_3')
// (5, 5, 'neigh_op_top_3')
// (5, 6, 'lutff_3/out')
// (5, 7, 'local_g0_3')
// (5, 7, 'lutff_1/in_2')
// (5, 7, 'neigh_op_bot_3')
// (6, 5, 'neigh_op_tnl_3')
// (6, 6, 'neigh_op_lft_3')
// (6, 7, 'neigh_op_bnl_3')

wire n182;
// (4, 5, 'neigh_op_tnr_4')
// (4, 6, 'neigh_op_rgt_4')
// (4, 7, 'neigh_op_bnr_4')
// (5, 5, 'local_g1_4')
// (5, 5, 'lutff_0/in_3')
// (5, 5, 'neigh_op_top_4')
// (5, 6, 'lutff_4/out')
// (5, 7, 'neigh_op_bot_4')
// (6, 5, 'neigh_op_tnl_4')
// (6, 6, 'neigh_op_lft_4')
// (6, 7, 'neigh_op_bnl_4')

wire n183;
// (4, 5, 'neigh_op_tnr_5')
// (4, 5, 'sp4_r_v_b_39')
// (4, 6, 'neigh_op_rgt_5')
// (4, 6, 'sp4_r_v_b_26')
// (4, 7, 'neigh_op_bnr_5')
// (4, 7, 'sp4_r_v_b_15')
// (4, 8, 'sp4_r_v_b_2')
// (5, 4, 'sp4_v_t_39')
// (5, 5, 'neigh_op_top_5')
// (5, 5, 'sp4_v_b_39')
// (5, 6, 'lutff_5/out')
// (5, 6, 'sp4_v_b_26')
// (5, 7, 'local_g1_5')
// (5, 7, 'lutff_1/in_1')
// (5, 7, 'neigh_op_bot_5')
// (5, 7, 'sp4_v_b_15')
// (5, 8, 'local_g0_2')
// (5, 8, 'lutff_0/in_2')
// (5, 8, 'lutff_4/in_2')
// (5, 8, 'sp4_v_b_2')
// (6, 5, 'neigh_op_tnl_5')
// (6, 6, 'neigh_op_lft_5')
// (6, 7, 'neigh_op_bnl_5')

wire n184;
// (4, 5, 'sp4_h_r_6')
// (5, 5, 'local_g0_3')
// (5, 5, 'local_g1_3')
// (5, 5, 'lutff_1/in_3')
// (5, 5, 'lutff_6/in_1')
// (5, 5, 'sp4_h_r_19')
// (6, 5, 'neigh_op_tnr_5')
// (6, 5, 'sp4_h_r_30')
// (6, 6, 'neigh_op_rgt_5')
// (6, 7, 'neigh_op_bnr_5')
// (7, 5, 'local_g1_5')
// (7, 5, 'lutff_1/in_3')
// (7, 5, 'lutff_4/in_0')
// (7, 5, 'neigh_op_top_5')
// (7, 5, 'sp4_h_r_43')
// (7, 6, 'lutff_5/out')
// (7, 6, 'sp4_r_v_b_43')
// (7, 7, 'neigh_op_bot_5')
// (7, 7, 'sp4_r_v_b_30')
// (7, 8, 'sp4_r_v_b_19')
// (7, 9, 'sp4_r_v_b_6')
// (8, 5, 'neigh_op_tnl_5')
// (8, 5, 'sp4_h_l_43')
// (8, 5, 'sp4_v_t_43')
// (8, 6, 'neigh_op_lft_5')
// (8, 6, 'sp4_v_b_43')
// (8, 7, 'neigh_op_bnl_5')
// (8, 7, 'sp4_v_b_30')
// (8, 8, 'sp4_v_b_19')
// (8, 9, 'sp4_v_b_6')

wire n185;
// (4, 5, 'sp4_h_r_8')
// (5, 5, 'sp4_h_r_21')
// (6, 5, 'sp4_h_r_32')
// (7, 2, 'sp4_r_v_b_39')
// (7, 3, 'local_g1_2')
// (7, 3, 'lutff_2/in_1')
// (7, 3, 'sp4_r_v_b_26')
// (7, 4, 'sp4_r_v_b_15')
// (7, 5, 'sp4_h_r_45')
// (7, 5, 'sp4_r_v_b_2')
// (8, 1, 'sp4_v_t_39')
// (8, 2, 'sp4_v_b_39')
// (8, 3, 'sp4_v_b_26')
// (8, 4, 'sp4_v_b_15')
// (8, 5, 'sp4_h_l_45')
// (8, 5, 'sp4_h_r_8')
// (8, 5, 'sp4_v_b_2')
// (9, 5, 'local_g0_5')
// (9, 5, 'lutff_1/in_0')
// (9, 5, 'sp4_h_r_21')
// (10, 3, 'neigh_op_tnr_2')
// (10, 4, 'neigh_op_rgt_2')
// (10, 5, 'neigh_op_bnr_2')
// (10, 5, 'sp4_h_r_32')
// (11, 2, 'sp4_r_v_b_45')
// (11, 3, 'neigh_op_top_2')
// (11, 3, 'sp4_r_v_b_32')
// (11, 4, 'local_g2_2')
// (11, 4, 'lutff_1/in_1')
// (11, 4, 'lutff_2/out')
// (11, 4, 'sp4_r_v_b_21')
// (11, 5, 'local_g0_2')
// (11, 5, 'lutff_1/in_1')
// (11, 5, 'neigh_op_bot_2')
// (11, 5, 'sp4_h_r_45')
// (11, 5, 'sp4_r_v_b_8')
// (12, 1, 'sp4_v_t_45')
// (12, 2, 'sp4_v_b_45')
// (12, 3, 'neigh_op_tnl_2')
// (12, 3, 'sp4_v_b_32')
// (12, 4, 'neigh_op_lft_2')
// (12, 4, 'sp4_v_b_21')
// (12, 5, 'neigh_op_bnl_2')
// (12, 5, 'sp4_h_l_45')
// (12, 5, 'sp4_v_b_8')

reg n186 = 0;
// (4, 6, 'local_g3_5')
// (4, 6, 'lutff_2/in_0')
// (4, 6, 'neigh_op_tnr_5')
// (4, 7, 'neigh_op_rgt_5')
// (4, 8, 'neigh_op_bnr_5')
// (5, 6, 'neigh_op_top_5')
// (5, 7, 'lutff_5/out')
// (5, 8, 'neigh_op_bot_5')
// (6, 6, 'neigh_op_tnl_5')
// (6, 7, 'neigh_op_lft_5')
// (6, 8, 'neigh_op_bnl_5')

wire n187;
// (4, 6, 'neigh_op_tnr_0')
// (4, 6, 'sp4_r_v_b_45')
// (4, 7, 'neigh_op_rgt_0')
// (4, 7, 'sp4_r_v_b_32')
// (4, 8, 'neigh_op_bnr_0')
// (4, 8, 'sp4_r_v_b_21')
// (4, 9, 'local_g2_0')
// (4, 9, 'lutff_2/in_2')
// (4, 9, 'sp4_r_v_b_8')
// (5, 5, 'sp4_v_t_45')
// (5, 6, 'neigh_op_top_0')
// (5, 6, 'sp4_v_b_45')
// (5, 7, 'lutff_0/out')
// (5, 7, 'sp4_v_b_32')
// (5, 8, 'local_g1_0')
// (5, 8, 'lutff_0/in_1')
// (5, 8, 'neigh_op_bot_0')
// (5, 8, 'sp4_v_b_21')
// (5, 9, 'sp4_v_b_8')
// (6, 6, 'neigh_op_tnl_0')
// (6, 7, 'neigh_op_lft_0')
// (6, 8, 'neigh_op_bnl_0')

wire n188;
// (4, 6, 'neigh_op_tnr_1')
// (4, 7, 'neigh_op_rgt_1')
// (4, 8, 'neigh_op_bnr_1')
// (5, 5, 'sp4_r_v_b_43')
// (5, 6, 'neigh_op_top_1')
// (5, 6, 'sp4_r_v_b_30')
// (5, 6, 'sp4_r_v_b_46')
// (5, 7, 'lutff_1/out')
// (5, 7, 'sp4_r_v_b_19')
// (5, 7, 'sp4_r_v_b_35')
// (5, 8, 'neigh_op_bot_1')
// (5, 8, 'sp4_r_v_b_22')
// (5, 8, 'sp4_r_v_b_6')
// (5, 9, 'sp4_r_v_b_11')
// (6, 4, 'sp4_v_t_43')
// (6, 5, 'sp4_v_b_43')
// (6, 5, 'sp4_v_t_46')
// (6, 6, 'neigh_op_tnl_1')
// (6, 6, 'sp4_v_b_30')
// (6, 6, 'sp4_v_b_46')
// (6, 7, 'neigh_op_lft_1')
// (6, 7, 'sp4_v_b_19')
// (6, 7, 'sp4_v_b_35')
// (6, 8, 'neigh_op_bnl_1')
// (6, 8, 'sp4_h_r_6')
// (6, 8, 'sp4_v_b_22')
// (6, 8, 'sp4_v_b_6')
// (6, 9, 'local_g0_3')
// (6, 9, 'local_g1_3')
// (6, 9, 'lutff_5/in_2')
// (6, 9, 'lutff_6/in_3')
// (6, 9, 'lutff_7/in_3')
// (6, 9, 'sp4_h_r_5')
// (6, 9, 'sp4_v_b_11')
// (7, 8, 'local_g0_3')
// (7, 8, 'local_g1_3')
// (7, 8, 'lutff_2/in_2')
// (7, 8, 'lutff_6/in_3')
// (7, 8, 'sp4_h_r_19')
// (7, 9, 'sp4_h_r_16')
// (8, 8, 'sp4_h_r_30')
// (8, 9, 'sp4_h_r_29')
// (9, 8, 'sp4_h_r_43')
// (9, 9, 'sp4_h_r_40')
// (10, 8, 'sp4_h_l_43')
// (10, 9, 'sp4_h_l_40')
// (10, 9, 'sp4_h_r_5')
// (11, 9, 'local_g0_0')
// (11, 9, 'lutff_4/in_2')
// (11, 9, 'sp4_h_r_16')
// (12, 9, 'sp4_h_r_29')
// (13, 9, 'span4_horz_29')

reg n189 = 0;
// (4, 6, 'neigh_op_tnr_2')
// (4, 7, 'neigh_op_rgt_2')
// (4, 8, 'neigh_op_bnr_2')
// (5, 6, 'neigh_op_top_2')
// (5, 7, 'lutff_2/out')
// (5, 7, 'sp4_h_r_4')
// (5, 8, 'neigh_op_bot_2')
// (6, 6, 'neigh_op_tnl_2')
// (6, 7, 'local_g1_1')
// (6, 7, 'lutff_6/in_0')
// (6, 7, 'neigh_op_lft_2')
// (6, 7, 'sp4_h_r_17')
// (6, 8, 'neigh_op_bnl_2')
// (7, 7, 'sp4_h_r_28')
// (8, 7, 'sp4_h_r_41')
// (9, 7, 'sp4_h_l_41')

reg n190 = 0;
// (4, 6, 'neigh_op_tnr_3')
// (4, 7, 'neigh_op_rgt_3')
// (4, 8, 'neigh_op_bnr_3')
// (5, 6, 'neigh_op_top_3')
// (5, 7, 'local_g2_3')
// (5, 7, 'lutff_3/out')
// (5, 7, 'lutff_7/in_0')
// (5, 8, 'neigh_op_bot_3')
// (6, 6, 'neigh_op_tnl_3')
// (6, 7, 'neigh_op_lft_3')
// (6, 8, 'neigh_op_bnl_3')

reg n191 = 0;
// (4, 6, 'neigh_op_tnr_7')
// (4, 7, 'neigh_op_rgt_7')
// (4, 8, 'neigh_op_bnr_7')
// (5, 6, 'neigh_op_top_7')
// (5, 7, 'local_g2_7')
// (5, 7, 'lutff_4/in_1')
// (5, 7, 'lutff_7/out')
// (5, 8, 'neigh_op_bot_7')
// (6, 6, 'neigh_op_tnl_7')
// (6, 7, 'local_g1_7')
// (6, 7, 'lutff_1/in_1')
// (6, 7, 'neigh_op_lft_7')
// (6, 8, 'neigh_op_bnl_7')

wire n192;
// (4, 6, 'sp4_r_v_b_38')
// (4, 7, 'sp4_r_v_b_27')
// (4, 8, 'sp4_r_v_b_14')
// (4, 9, 'sp4_r_v_b_3')
// (4, 10, 'sp4_r_v_b_42')
// (4, 11, 'neigh_op_tnr_1')
// (4, 11, 'sp4_r_v_b_31')
// (4, 12, 'neigh_op_rgt_1')
// (4, 12, 'sp4_r_v_b_18')
// (4, 13, 'neigh_op_bnr_1')
// (4, 13, 'sp4_r_v_b_7')
// (5, 5, 'sp4_v_t_38')
// (5, 6, 'sp4_v_b_38')
// (5, 7, 'sp4_v_b_27')
// (5, 8, 'sp4_v_b_14')
// (5, 9, 'local_g0_3')
// (5, 9, 'lutff_0/in_3')
// (5, 9, 'sp4_v_b_3')
// (5, 9, 'sp4_v_t_42')
// (5, 10, 'sp4_v_b_42')
// (5, 11, 'neigh_op_top_1')
// (5, 11, 'sp4_v_b_31')
// (5, 12, 'lutff_1/out')
// (5, 12, 'sp4_v_b_18')
// (5, 13, 'neigh_op_bot_1')
// (5, 13, 'sp4_v_b_7')
// (6, 11, 'neigh_op_tnl_1')
// (6, 12, 'neigh_op_lft_1')
// (6, 13, 'neigh_op_bnl_1')

wire n193;
// (4, 6, 'sp4_r_v_b_40')
// (4, 7, 'neigh_op_tnr_0')
// (4, 7, 'sp4_r_v_b_29')
// (4, 8, 'local_g3_0')
// (4, 8, 'lutff_2/in_3')
// (4, 8, 'lutff_4/in_3')
// (4, 8, 'neigh_op_rgt_0')
// (4, 8, 'sp4_r_v_b_16')
// (4, 9, 'local_g1_0')
// (4, 9, 'local_g1_5')
// (4, 9, 'lutff_1/in_3')
// (4, 9, 'lutff_7/in_2')
// (4, 9, 'neigh_op_bnr_0')
// (4, 9, 'sp4_r_v_b_5')
// (5, 5, 'sp4_v_t_40')
// (5, 6, 'sp4_v_b_40')
// (5, 7, 'neigh_op_top_0')
// (5, 7, 'sp4_r_v_b_44')
// (5, 7, 'sp4_v_b_29')
// (5, 8, 'lutff_0/out')
// (5, 8, 'sp4_r_v_b_33')
// (5, 8, 'sp4_v_b_16')
// (5, 9, 'neigh_op_bot_0')
// (5, 9, 'sp4_r_v_b_20')
// (5, 9, 'sp4_v_b_5')
// (5, 10, 'sp4_r_v_b_9')
// (6, 6, 'sp4_v_t_44')
// (6, 7, 'neigh_op_tnl_0')
// (6, 7, 'sp4_v_b_44')
// (6, 8, 'neigh_op_lft_0')
// (6, 8, 'sp4_v_b_33')
// (6, 9, 'neigh_op_bnl_0')
// (6, 9, 'sp4_v_b_20')
// (6, 10, 'sp4_h_r_9')
// (6, 10, 'sp4_v_b_9')
// (7, 10, 'local_g0_4')
// (7, 10, 'lutff_7/in_3')
// (7, 10, 'sp4_h_r_20')
// (8, 10, 'sp4_h_r_33')
// (9, 10, 'sp4_h_r_44')
// (10, 10, 'sp4_h_l_44')

wire n194;
// (4, 7, 'neigh_op_tnr_3')
// (4, 8, 'local_g3_3')
// (4, 8, 'lutff_2/in_2')
// (4, 8, 'lutff_3/in_3')
// (4, 8, 'neigh_op_rgt_3')
// (4, 9, 'neigh_op_bnr_3')
// (5, 7, 'neigh_op_top_3')
// (5, 8, 'lutff_3/out')
// (5, 9, 'neigh_op_bot_3')
// (6, 7, 'neigh_op_tnl_3')
// (6, 8, 'neigh_op_lft_3')
// (6, 9, 'neigh_op_bnl_3')

wire n195;
// (4, 7, 'neigh_op_tnr_4')
// (4, 8, 'local_g2_4')
// (4, 8, 'lutff_1/in_3')
// (4, 8, 'lutff_6/in_2')
// (4, 8, 'neigh_op_rgt_4')
// (4, 9, 'local_g0_4')
// (4, 9, 'lutff_3/in_3')
// (4, 9, 'lutff_5/in_3')
// (4, 9, 'neigh_op_bnr_4')
// (5, 7, 'neigh_op_top_4')
// (5, 8, 'lutff_4/out')
// (5, 9, 'local_g0_4')
// (5, 9, 'lutff_3/in_3')
// (5, 9, 'neigh_op_bot_4')
// (6, 7, 'neigh_op_tnl_4')
// (6, 8, 'neigh_op_lft_4')
// (6, 9, 'neigh_op_bnl_4')

reg n196 = 0;
// (4, 7, 'neigh_op_tnr_6')
// (4, 8, 'neigh_op_rgt_6')
// (4, 9, 'neigh_op_bnr_6')
// (5, 7, 'local_g1_6')
// (5, 7, 'lutff_5/in_0')
// (5, 7, 'neigh_op_top_6')
// (5, 8, 'lutff_6/out')
// (5, 9, 'neigh_op_bot_6')
// (6, 7, 'neigh_op_tnl_6')
// (6, 8, 'neigh_op_lft_6')
// (6, 9, 'neigh_op_bnl_6')

reg n197 = 0;
// (4, 7, 'neigh_op_tnr_7')
// (4, 8, 'neigh_op_rgt_7')
// (4, 9, 'neigh_op_bnr_7')
// (5, 3, 'sp12_v_t_22')
// (5, 4, 'sp12_v_b_22')
// (5, 5, 'sp12_v_b_21')
// (5, 6, 'sp12_v_b_18')
// (5, 7, 'local_g3_1')
// (5, 7, 'lutff_6/in_0')
// (5, 7, 'neigh_op_top_7')
// (5, 7, 'sp12_v_b_17')
// (5, 8, 'lutff_7/out')
// (5, 8, 'sp12_v_b_14')
// (5, 9, 'neigh_op_bot_7')
// (5, 9, 'sp12_v_b_13')
// (5, 10, 'sp12_v_b_10')
// (5, 11, 'sp12_v_b_9')
// (5, 12, 'sp12_v_b_6')
// (5, 13, 'sp12_v_b_5')
// (5, 14, 'sp12_v_b_2')
// (5, 15, 'sp12_v_b_1')
// (6, 7, 'neigh_op_tnl_7')
// (6, 8, 'neigh_op_lft_7')
// (6, 9, 'neigh_op_bnl_7')

reg n198 = 0;
// (4, 7, 'sp12_h_r_0')
// (5, 6, 'neigh_op_tnr_6')
// (5, 7, 'neigh_op_rgt_6')
// (5, 7, 'sp12_h_r_3')
// (5, 8, 'neigh_op_bnr_6')
// (6, 5, 'sp4_r_v_b_37')
// (6, 6, 'neigh_op_top_6')
// (6, 6, 'sp4_r_v_b_24')
// (6, 7, 'lutff_6/out')
// (6, 7, 'sp12_h_r_4')
// (6, 7, 'sp4_r_v_b_13')
// (6, 8, 'neigh_op_bot_6')
// (6, 8, 'sp4_r_v_b_0')
// (7, 4, 'sp4_v_t_37')
// (7, 5, 'sp4_v_b_37')
// (7, 6, 'neigh_op_tnl_6')
// (7, 6, 'sp4_v_b_24')
// (7, 7, 'local_g0_5')
// (7, 7, 'lutff_7/in_0')
// (7, 7, 'neigh_op_lft_6')
// (7, 7, 'sp12_h_r_7')
// (7, 7, 'sp4_v_b_13')
// (7, 8, 'neigh_op_bnl_6')
// (7, 8, 'sp4_v_b_0')
// (8, 7, 'local_g1_0')
// (8, 7, 'lutff_4/in_3')
// (8, 7, 'sp12_h_r_8')
// (9, 7, 'sp12_h_r_11')
// (10, 7, 'sp12_h_r_12')
// (11, 7, 'sp12_h_r_15')
// (12, 7, 'sp12_h_r_16')
// (13, 7, 'span12_horz_16')

reg n199 = 0;
// (4, 7, 'sp4_h_r_7')
// (5, 7, 'local_g0_2')
// (5, 7, 'lutff_4/in_0')
// (5, 7, 'sp4_h_r_18')
// (6, 6, 'neigh_op_tnr_5')
// (6, 7, 'local_g2_7')
// (6, 7, 'local_g3_7')
// (6, 7, 'lutff_4/in_0')
// (6, 7, 'lutff_7/in_0')
// (6, 7, 'neigh_op_rgt_5')
// (6, 7, 'sp4_h_r_31')
// (6, 8, 'neigh_op_bnr_5')
// (7, 6, 'neigh_op_top_5')
// (7, 7, 'local_g1_5')
// (7, 7, 'lutff_5/out')
// (7, 7, 'lutff_6/in_0')
// (7, 7, 'sp4_h_r_42')
// (7, 8, 'neigh_op_bot_5')
// (8, 6, 'neigh_op_tnl_5')
// (8, 7, 'neigh_op_lft_5')
// (8, 7, 'sp4_h_l_42')
// (8, 8, 'neigh_op_bnl_5')

wire n200;
// (4, 8, 'neigh_op_tnr_1')
// (4, 9, 'neigh_op_rgt_1')
// (4, 10, 'neigh_op_bnr_1')
// (5, 6, 'sp12_v_t_22')
// (5, 7, 'sp12_v_b_22')
// (5, 8, 'neigh_op_top_1')
// (5, 8, 'sp12_v_b_21')
// (5, 9, 'lutff_1/out')
// (5, 9, 'sp12_v_b_18')
// (5, 10, 'neigh_op_bot_1')
// (5, 10, 'sp12_v_b_17')
// (5, 11, 'local_g2_6')
// (5, 11, 'lutff_3/in_3')
// (5, 11, 'sp12_v_b_14')
// (5, 12, 'sp12_v_b_13')
// (5, 13, 'sp12_v_b_10')
// (5, 14, 'sp12_v_b_9')
// (5, 15, 'sp12_v_b_6')
// (5, 16, 'sp12_v_b_5')
// (5, 17, 'span12_vert_2')
// (6, 8, 'neigh_op_tnl_1')
// (6, 9, 'local_g1_1')
// (6, 9, 'lutff_3/in_3')
// (6, 9, 'lutff_5/in_3')
// (6, 9, 'neigh_op_lft_1')
// (6, 10, 'neigh_op_bnl_1')

reg \d_out[4] = 0 ;
// (4, 8, 'neigh_op_tnr_3')
// (4, 9, 'neigh_op_rgt_3')
// (4, 10, 'neigh_op_bnr_3')
// (5, 8, 'neigh_op_top_3')
// (5, 9, 'lutff_3/out')
// (5, 9, 'sp4_h_r_6')
// (5, 10, 'neigh_op_bot_3')
// (6, 8, 'neigh_op_tnl_3')
// (6, 9, 'neigh_op_lft_3')
// (6, 9, 'sp4_h_r_19')
// (6, 10, 'neigh_op_bnl_3')
// (7, 9, 'sp4_h_r_30')
// (8, 9, 'sp4_h_r_43')
// (9, 9, 'sp4_h_l_43')
// (9, 9, 'sp4_h_r_6')
// (10, 9, 'sp4_h_r_19')
// (11, 9, 'sp4_h_r_30')
// (12, 9, 'sp4_h_r_43')
// (13, 9, 'io_1/D_OUT_0')
// (13, 9, 'io_1/PAD')
// (13, 9, 'local_g0_3')
// (13, 9, 'span4_horz_43')

reg n202 = 0;
// (4, 8, 'neigh_op_tnr_4')
// (4, 9, 'neigh_op_rgt_4')
// (4, 10, 'neigh_op_bnr_4')
// (5, 8, 'neigh_op_top_4')
// (5, 9, 'local_g2_4')
// (5, 9, 'lutff_4/out')
// (5, 9, 'lutff_6/in_0')
// (5, 10, 'neigh_op_bot_4')
// (6, 8, 'neigh_op_tnl_4')
// (6, 9, 'neigh_op_lft_4')
// (6, 10, 'neigh_op_bnl_4')

reg n203 = 0;
// (4, 8, 'neigh_op_tnr_5')
// (4, 9, 'neigh_op_rgt_5')
// (4, 10, 'neigh_op_bnr_5')
// (5, 8, 'local_g1_5')
// (5, 8, 'lutff_6/in_0')
// (5, 8, 'neigh_op_top_5')
// (5, 9, 'lutff_5/out')
// (5, 10, 'neigh_op_bot_5')
// (6, 8, 'neigh_op_tnl_5')
// (6, 9, 'neigh_op_lft_5')
// (6, 10, 'neigh_op_bnl_5')

reg n204 = 0;
// (4, 8, 'neigh_op_tnr_6')
// (4, 9, 'neigh_op_rgt_6')
// (4, 10, 'neigh_op_bnr_6')
// (5, 8, 'local_g1_6')
// (5, 8, 'lutff_7/in_0')
// (5, 8, 'neigh_op_top_6')
// (5, 9, 'lutff_6/out')
// (5, 10, 'neigh_op_bot_6')
// (6, 8, 'neigh_op_tnl_6')
// (6, 9, 'neigh_op_lft_6')
// (6, 10, 'neigh_op_bnl_6')

reg n205 = 0;
// (4, 9, 'neigh_op_tnr_0')
// (4, 10, 'neigh_op_rgt_0')
// (4, 11, 'neigh_op_bnr_0')
// (5, 9, 'neigh_op_top_0')
// (5, 10, 'local_g1_0')
// (5, 10, 'lutff_0/out')
// (5, 10, 'lutff_7/in_0')
// (5, 11, 'neigh_op_bot_0')
// (6, 9, 'neigh_op_tnl_0')
// (6, 10, 'neigh_op_lft_0')
// (6, 11, 'neigh_op_bnl_0')

reg n206 = 0;
// (4, 9, 'neigh_op_tnr_1')
// (4, 10, 'neigh_op_rgt_1')
// (4, 11, 'neigh_op_bnr_1')
// (5, 9, 'neigh_op_top_1')
// (5, 10, 'local_g3_1')
// (5, 10, 'lutff_0/in_0')
// (5, 10, 'lutff_1/out')
// (5, 11, 'neigh_op_bot_1')
// (6, 9, 'neigh_op_tnl_1')
// (6, 10, 'neigh_op_lft_1')
// (6, 11, 'neigh_op_bnl_1')

reg n207 = 0;
// (4, 9, 'neigh_op_tnr_2')
// (4, 10, 'neigh_op_rgt_2')
// (4, 11, 'neigh_op_bnr_2')
// (5, 9, 'neigh_op_top_2')
// (5, 10, 'local_g0_2')
// (5, 10, 'lutff_2/out')
// (5, 10, 'lutff_6/in_0')
// (5, 11, 'neigh_op_bot_2')
// (6, 9, 'neigh_op_tnl_2')
// (6, 10, 'neigh_op_lft_2')
// (6, 11, 'neigh_op_bnl_2')

reg n208 = 0;
// (4, 9, 'neigh_op_tnr_3')
// (4, 10, 'neigh_op_rgt_3')
// (4, 11, 'neigh_op_bnr_3')
// (5, 9, 'neigh_op_top_3')
// (5, 10, 'local_g1_3')
// (5, 10, 'lutff_2/in_0')
// (5, 10, 'lutff_3/out')
// (5, 11, 'neigh_op_bot_3')
// (6, 9, 'neigh_op_tnl_3')
// (6, 10, 'neigh_op_lft_3')
// (6, 11, 'neigh_op_bnl_3')

reg n209 = 0;
// (4, 9, 'neigh_op_tnr_5')
// (4, 10, 'neigh_op_rgt_5')
// (4, 11, 'neigh_op_bnr_5')
// (5, 9, 'local_g0_5')
// (5, 9, 'lutff_2/in_3')
// (5, 9, 'neigh_op_top_5')
// (5, 10, 'lutff_5/out')
// (5, 11, 'neigh_op_bot_5')
// (6, 9, 'neigh_op_tnl_5')
// (6, 10, 'neigh_op_lft_5')
// (6, 11, 'neigh_op_bnl_5')

reg n210 = 0;
// (4, 9, 'neigh_op_tnr_6')
// (4, 10, 'neigh_op_rgt_6')
// (4, 11, 'neigh_op_bnr_6')
// (5, 9, 'neigh_op_top_6')
// (5, 10, 'lutff_6/out')
// (5, 11, 'local_g1_6')
// (5, 11, 'lutff_5/in_0')
// (5, 11, 'neigh_op_bot_6')
// (6, 9, 'neigh_op_tnl_6')
// (6, 10, 'neigh_op_lft_6')
// (6, 11, 'neigh_op_bnl_6')

reg n211 = 0;
// (4, 9, 'neigh_op_tnr_7')
// (4, 10, 'neigh_op_rgt_7')
// (4, 11, 'neigh_op_bnr_7')
// (5, 9, 'neigh_op_top_7')
// (5, 10, 'local_g0_7')
// (5, 10, 'lutff_5/in_0')
// (5, 10, 'lutff_7/out')
// (5, 11, 'neigh_op_bot_7')
// (6, 9, 'neigh_op_tnl_7')
// (6, 10, 'neigh_op_lft_7')
// (6, 11, 'neigh_op_bnl_7')

reg n212 = 0;
// (4, 9, 'sp12_h_r_1')
// (5, 9, 'sp12_h_r_2')
// (6, 9, 'sp12_h_r_5')
// (7, 9, 'local_g1_6')
// (7, 9, 'lutff_7/in_0')
// (7, 9, 'sp12_h_r_6')
// (8, 9, 'sp12_h_r_9')
// (9, 9, 'sp12_h_r_10')
// (10, 8, 'neigh_op_tnr_3')
// (10, 9, 'neigh_op_rgt_3')
// (10, 9, 'sp12_h_r_13')
// (10, 10, 'neigh_op_bnr_3')
// (11, 8, 'neigh_op_top_3')
// (11, 9, 'lutff_3/out')
// (11, 9, 'sp12_h_r_14')
// (11, 10, 'neigh_op_bot_3')
// (12, 8, 'neigh_op_tnl_3')
// (12, 9, 'neigh_op_lft_3')
// (12, 9, 'sp12_h_r_17')
// (12, 10, 'neigh_op_bnl_3')
// (13, 9, 'span12_horz_17')

reg n213 = 0;
// (4, 9, 'sp4_h_r_2')
// (5, 9, 'local_g1_7')
// (5, 9, 'lutff_4/in_0')
// (5, 9, 'sp4_h_r_15')
// (6, 8, 'neigh_op_tnr_4')
// (6, 9, 'neigh_op_rgt_4')
// (6, 9, 'sp4_h_r_26')
// (6, 10, 'neigh_op_bnr_4')
// (7, 6, 'sp4_r_v_b_44')
// (7, 7, 'sp4_r_v_b_33')
// (7, 8, 'neigh_op_top_4')
// (7, 8, 'sp4_r_v_b_20')
// (7, 9, 'lutff_4/out')
// (7, 9, 'sp4_h_r_39')
// (7, 9, 'sp4_r_v_b_9')
// (7, 10, 'neigh_op_bot_4')
// (8, 5, 'sp4_v_t_44')
// (8, 6, 'sp4_v_b_44')
// (8, 7, 'sp4_v_b_33')
// (8, 8, 'neigh_op_tnl_4')
// (8, 8, 'sp4_v_b_20')
// (8, 9, 'neigh_op_lft_4')
// (8, 9, 'sp4_h_l_39')
// (8, 9, 'sp4_v_b_9')
// (8, 10, 'neigh_op_bnl_4')

wire n214;
// (4, 10, 'neigh_op_tnr_0')
// (4, 11, 'neigh_op_rgt_0')
// (4, 12, 'neigh_op_bnr_0')
// (5, 10, 'neigh_op_top_0')
// (5, 11, 'lutff_0/out')
// (5, 12, 'local_g0_0')
// (5, 12, 'local_g1_0')
// (5, 12, 'lutff_4/in_1')
// (5, 12, 'lutff_5/in_1')
// (5, 12, 'neigh_op_bot_0')
// (6, 10, 'neigh_op_tnl_0')
// (6, 11, 'neigh_op_lft_0')
// (6, 12, 'neigh_op_bnl_0')

reg n215 = 0;
// (4, 10, 'neigh_op_tnr_2')
// (4, 11, 'neigh_op_rgt_2')
// (4, 12, 'neigh_op_bnr_2')
// (5, 10, 'neigh_op_top_2')
// (5, 11, 'local_g0_2')
// (5, 11, 'local_g1_2')
// (5, 11, 'lutff_2/out')
// (5, 11, 'lutff_4/in_2')
// (5, 11, 'lutff_6/in_1')
// (5, 12, 'neigh_op_bot_2')
// (6, 10, 'neigh_op_tnl_2')
// (6, 11, 'neigh_op_lft_2')
// (6, 12, 'neigh_op_bnl_2')

reg n216 = 0;
// (4, 10, 'neigh_op_tnr_3')
// (4, 11, 'neigh_op_rgt_3')
// (4, 12, 'neigh_op_bnr_3')
// (5, 10, 'neigh_op_top_3')
// (5, 11, 'local_g0_3')
// (5, 11, 'lutff_2/in_1')
// (5, 11, 'lutff_3/out')
// (5, 11, 'lutff_7/in_2')
// (5, 12, 'neigh_op_bot_3')
// (6, 10, 'neigh_op_tnl_3')
// (6, 11, 'neigh_op_lft_3')
// (6, 12, 'neigh_op_bnl_3')

reg n217 = 0;
// (4, 10, 'neigh_op_tnr_4')
// (4, 11, 'neigh_op_rgt_4')
// (4, 12, 'neigh_op_bnr_4')
// (5, 10, 'neigh_op_top_4')
// (5, 11, 'local_g1_4')
// (5, 11, 'lutff_0/in_1')
// (5, 11, 'lutff_4/out')
// (5, 12, 'neigh_op_bot_4')
// (6, 10, 'neigh_op_tnl_4')
// (6, 11, 'neigh_op_lft_4')
// (6, 12, 'neigh_op_bnl_4')

reg n218 = 0;
// (4, 10, 'neigh_op_tnr_5')
// (4, 10, 'sp4_r_v_b_39')
// (4, 11, 'neigh_op_rgt_5')
// (4, 11, 'sp4_r_v_b_26')
// (4, 11, 'sp4_r_v_b_42')
// (4, 12, 'neigh_op_bnr_5')
// (4, 12, 'sp4_r_v_b_15')
// (4, 12, 'sp4_r_v_b_31')
// (4, 13, 'sp4_r_v_b_18')
// (4, 13, 'sp4_r_v_b_2')
// (4, 14, 'sp4_r_v_b_7')
// (5, 9, 'sp4_v_t_39')
// (5, 10, 'neigh_op_top_5')
// (5, 10, 'sp4_v_b_39')
// (5, 10, 'sp4_v_t_42')
// (5, 11, 'lutff_5/out')
// (5, 11, 'sp4_v_b_26')
// (5, 11, 'sp4_v_b_42')
// (5, 12, 'local_g0_7')
// (5, 12, 'lutff_0/in_1')
// (5, 12, 'neigh_op_bot_5')
// (5, 12, 'sp4_v_b_15')
// (5, 12, 'sp4_v_b_31')
// (5, 13, 'sp4_v_b_18')
// (5, 13, 'sp4_v_b_2')
// (5, 14, 'local_g1_7')
// (5, 14, 'lutff_5/in_1')
// (5, 14, 'sp4_v_b_7')
// (6, 10, 'neigh_op_tnl_5')
// (6, 11, 'neigh_op_lft_5')
// (6, 12, 'neigh_op_bnl_5')

reg n219 = 0;
// (4, 10, 'neigh_op_tnr_6')
// (4, 11, 'neigh_op_rgt_6')
// (4, 12, 'neigh_op_bnr_6')
// (5, 10, 'neigh_op_top_6')
// (5, 11, 'local_g0_6')
// (5, 11, 'lutff_0/in_2')
// (5, 11, 'lutff_1/in_1')
// (5, 11, 'lutff_6/out')
// (5, 12, 'neigh_op_bot_6')
// (6, 10, 'neigh_op_tnl_6')
// (6, 11, 'neigh_op_lft_6')
// (6, 12, 'neigh_op_bnl_6')

reg n220 = 0;
// (4, 10, 'neigh_op_tnr_7')
// (4, 11, 'neigh_op_rgt_7')
// (4, 12, 'neigh_op_bnr_7')
// (5, 10, 'neigh_op_top_7')
// (5, 11, 'local_g0_7')
// (5, 11, 'lutff_4/in_1')
// (5, 11, 'lutff_7/out')
// (5, 12, 'neigh_op_bot_7')
// (6, 10, 'neigh_op_tnl_7')
// (6, 11, 'neigh_op_lft_7')
// (6, 12, 'neigh_op_bnl_7')

reg n221 = 0;
// (4, 10, 'sp4_r_v_b_45')
// (4, 11, 'sp4_r_v_b_32')
// (4, 12, 'sp4_r_v_b_21')
// (4, 13, 'sp4_r_v_b_8')
// (5, 9, 'local_g0_2')
// (5, 9, 'lutff_0/in_2')
// (5, 9, 'sp4_h_r_2')
// (5, 9, 'sp4_v_t_45')
// (5, 10, 'local_g2_5')
// (5, 10, 'lutff_3/in_2')
// (5, 10, 'sp4_v_b_45')
// (5, 11, 'sp4_v_b_32')
// (5, 12, 'sp4_v_b_21')
// (5, 13, 'sp4_v_b_8')
// (6, 9, 'sp4_h_r_15')
// (7, 9, 'sp4_h_r_26')
// (8, 5, 'local_g3_6')
// (8, 5, 'lutff_7/in_0')
// (8, 5, 'neigh_op_tnr_6')
// (8, 6, 'neigh_op_rgt_6')
// (8, 6, 'sp4_r_v_b_44')
// (8, 7, 'neigh_op_bnr_6')
// (8, 7, 'sp4_r_v_b_33')
// (8, 8, 'sp4_r_v_b_20')
// (8, 9, 'sp4_h_r_39')
// (8, 9, 'sp4_r_v_b_9')
// (8, 10, 'sp4_r_v_b_37')
// (8, 11, 'local_g0_0')
// (8, 11, 'lutff_4/in_0')
// (8, 11, 'sp4_r_v_b_24')
// (8, 12, 'sp4_r_v_b_13')
// (8, 13, 'sp4_r_v_b_0')
// (9, 5, 'neigh_op_top_6')
// (9, 5, 'sp4_v_t_44')
// (9, 6, 'lutff_6/out')
// (9, 6, 'sp4_v_b_44')
// (9, 7, 'neigh_op_bot_6')
// (9, 7, 'sp4_v_b_33')
// (9, 8, 'sp4_v_b_20')
// (9, 9, 'sp4_h_l_39')
// (9, 9, 'sp4_v_b_9')
// (9, 9, 'sp4_v_t_37')
// (9, 10, 'sp4_v_b_37')
// (9, 11, 'sp4_v_b_24')
// (9, 12, 'sp4_v_b_13')
// (9, 13, 'sp4_v_b_0')
// (10, 5, 'neigh_op_tnl_6')
// (10, 6, 'neigh_op_lft_6')
// (10, 7, 'neigh_op_bnl_6')

wire n222;
// (4, 11, 'neigh_op_tnr_0')
// (4, 12, 'neigh_op_rgt_0')
// (4, 13, 'neigh_op_bnr_0')
// (5, 11, 'neigh_op_top_0')
// (5, 12, 'local_g2_0')
// (5, 12, 'lutff_0/out')
// (5, 12, 'lutff_1/in_3')
// (5, 13, 'neigh_op_bot_0')
// (6, 11, 'neigh_op_tnl_0')
// (6, 12, 'neigh_op_lft_0')
// (6, 13, 'neigh_op_bnl_0')

wire n223;
// (4, 11, 'neigh_op_tnr_3')
// (4, 12, 'neigh_op_rgt_3')
// (4, 13, 'neigh_op_bnr_3')
// (5, 11, 'neigh_op_top_3')
// (5, 12, 'local_g0_3')
// (5, 12, 'lutff_3/out')
// (5, 12, 'lutff_4/in_3')
// (5, 13, 'neigh_op_bot_3')
// (6, 11, 'neigh_op_tnl_3')
// (6, 12, 'neigh_op_lft_3')
// (6, 13, 'neigh_op_bnl_3')

reg n224 = 0;
// (4, 11, 'neigh_op_tnr_5')
// (4, 12, 'neigh_op_rgt_5')
// (4, 13, 'neigh_op_bnr_5')
// (5, 11, 'neigh_op_top_5')
// (5, 12, 'local_g0_5')
// (5, 12, 'lutff_5/out')
// (5, 12, 'lutff_7/in_0')
// (5, 13, 'neigh_op_bot_5')
// (6, 11, 'neigh_op_tnl_5')
// (6, 12, 'neigh_op_lft_5')
// (6, 13, 'neigh_op_bnl_5')

reg n225 = 0;
// (4, 11, 'neigh_op_tnr_6')
// (4, 12, 'neigh_op_rgt_6')
// (4, 13, 'neigh_op_bnr_6')
// (5, 11, 'neigh_op_top_6')
// (5, 12, 'lutff_6/out')
// (5, 13, 'local_g0_6')
// (5, 13, 'lutff_4/in_0')
// (5, 13, 'neigh_op_bot_6')
// (6, 11, 'neigh_op_tnl_6')
// (6, 12, 'neigh_op_lft_6')
// (6, 13, 'neigh_op_bnl_6')

reg n226 = 0;
// (4, 11, 'neigh_op_tnr_7')
// (4, 12, 'neigh_op_rgt_7')
// (4, 13, 'neigh_op_bnr_7')
// (5, 11, 'neigh_op_top_7')
// (5, 12, 'local_g1_7')
// (5, 12, 'lutff_6/in_0')
// (5, 12, 'lutff_7/out')
// (5, 13, 'neigh_op_bot_7')
// (6, 11, 'neigh_op_tnl_7')
// (6, 12, 'neigh_op_lft_7')
// (6, 13, 'neigh_op_bnl_7')

reg n227 = 0;
// (4, 11, 'sp12_h_r_1')
// (5, 11, 'sp12_h_r_2')
// (6, 10, 'neigh_op_tnr_7')
// (6, 11, 'neigh_op_rgt_7')
// (6, 11, 'sp12_h_r_5')
// (6, 12, 'neigh_op_bnr_7')
// (7, 10, 'neigh_op_top_7')
// (7, 11, 'lutff_7/out')
// (7, 11, 'sp12_h_r_6')
// (7, 12, 'neigh_op_bot_7')
// (8, 10, 'neigh_op_tnl_7')
// (8, 11, 'neigh_op_lft_7')
// (8, 11, 'sp12_h_r_9')
// (8, 12, 'neigh_op_bnl_7')
// (9, 11, 'local_g1_2')
// (9, 11, 'lutff_1/in_2')
// (9, 11, 'sp12_h_r_10')
// (10, 11, 'sp12_h_r_13')
// (11, 11, 'sp12_h_r_14')
// (12, 11, 'sp12_h_r_17')
// (13, 11, 'span12_horz_17')

wire n228;
// (4, 12, 'neigh_op_tnr_0')
// (4, 13, 'neigh_op_rgt_0')
// (4, 14, 'neigh_op_bnr_0')
// (5, 11, 'sp4_r_v_b_41')
// (5, 12, 'local_g0_4')
// (5, 12, 'lutff_3/in_3')
// (5, 12, 'neigh_op_top_0')
// (5, 12, 'sp4_r_v_b_28')
// (5, 13, 'lutff_0/out')
// (5, 13, 'sp4_r_v_b_17')
// (5, 14, 'neigh_op_bot_0')
// (5, 14, 'sp4_r_v_b_4')
// (6, 10, 'sp4_v_t_41')
// (6, 11, 'sp4_v_b_41')
// (6, 12, 'neigh_op_tnl_0')
// (6, 12, 'sp4_v_b_28')
// (6, 13, 'neigh_op_lft_0')
// (6, 13, 'sp4_v_b_17')
// (6, 14, 'neigh_op_bnl_0')
// (6, 14, 'sp4_v_b_4')

reg n229 = 0;
// (4, 12, 'neigh_op_tnr_1')
// (4, 13, 'neigh_op_rgt_1')
// (4, 14, 'neigh_op_bnr_1')
// (5, 12, 'neigh_op_top_1')
// (5, 13, 'local_g3_1')
// (5, 13, 'lutff_1/out')
// (5, 13, 'lutff_6/in_0')
// (5, 14, 'neigh_op_bot_1')
// (6, 12, 'neigh_op_tnl_1')
// (6, 13, 'neigh_op_lft_1')
// (6, 14, 'neigh_op_bnl_1')

reg n230 = 0;
// (4, 12, 'neigh_op_tnr_2')
// (4, 13, 'neigh_op_rgt_2')
// (4, 14, 'neigh_op_bnr_2')
// (5, 12, 'neigh_op_top_2')
// (5, 13, 'local_g1_2')
// (5, 13, 'lutff_1/in_0')
// (5, 13, 'lutff_2/out')
// (5, 14, 'neigh_op_bot_2')
// (6, 12, 'neigh_op_tnl_2')
// (6, 13, 'neigh_op_lft_2')
// (6, 14, 'neigh_op_bnl_2')

reg n231 = 0;
// (4, 12, 'neigh_op_tnr_4')
// (4, 13, 'neigh_op_rgt_4')
// (4, 14, 'neigh_op_bnr_4')
// (5, 12, 'neigh_op_top_4')
// (5, 13, 'local_g1_4')
// (5, 13, 'lutff_0/in_1')
// (5, 13, 'lutff_2/in_1')
// (5, 13, 'lutff_4/out')
// (5, 14, 'neigh_op_bot_4')
// (6, 12, 'neigh_op_tnl_4')
// (6, 13, 'neigh_op_lft_4')
// (6, 14, 'neigh_op_bnl_4')

reg n232 = 0;
// (4, 12, 'neigh_op_tnr_6')
// (4, 13, 'neigh_op_rgt_6')
// (4, 14, 'neigh_op_bnr_6')
// (5, 12, 'neigh_op_top_6')
// (5, 13, 'local_g1_6')
// (5, 13, 'lutff_6/out')
// (5, 13, 'lutff_7/in_0')
// (5, 14, 'neigh_op_bot_6')
// (6, 12, 'neigh_op_tnl_6')
// (6, 13, 'neigh_op_lft_6')
// (6, 14, 'neigh_op_bnl_6')

reg n233 = 0;
// (4, 12, 'neigh_op_tnr_7')
// (4, 13, 'local_g3_7')
// (4, 13, 'lutff_5/in_1')
// (4, 13, 'neigh_op_rgt_7')
// (4, 14, 'neigh_op_bnr_7')
// (5, 12, 'neigh_op_top_7')
// (5, 13, 'local_g3_7')
// (5, 13, 'lutff_0/in_0')
// (5, 13, 'lutff_7/out')
// (5, 14, 'neigh_op_bot_7')
// (6, 12, 'neigh_op_tnl_7')
// (6, 13, 'neigh_op_lft_7')
// (6, 14, 'neigh_op_bnl_7')

reg n234 = 0;
// (4, 12, 'sp12_h_r_1')
// (5, 12, 'sp12_h_r_2')
// (6, 12, 'sp12_h_r_5')
// (7, 12, 'sp12_h_r_6')
// (8, 11, 'neigh_op_tnr_1')
// (8, 12, 'neigh_op_rgt_1')
// (8, 12, 'sp12_h_r_9')
// (8, 13, 'neigh_op_bnr_1')
// (9, 11, 'neigh_op_top_1')
// (9, 12, 'lutff_1/out')
// (9, 12, 'sp12_h_r_10')
// (9, 13, 'neigh_op_bot_1')
// (10, 11, 'neigh_op_tnl_1')
// (10, 12, 'neigh_op_lft_1')
// (10, 12, 'sp12_h_r_13')
// (10, 13, 'neigh_op_bnl_1')
// (11, 12, 'local_g1_6')
// (11, 12, 'lutff_7/in_0')
// (11, 12, 'sp12_h_r_14')
// (12, 12, 'sp12_h_r_17')
// (13, 12, 'span12_horz_17')

reg n235 = 0;
// (4, 13, 'neigh_op_tnr_2')
// (4, 14, 'local_g3_2')
// (4, 14, 'lutff_6/in_1')
// (4, 14, 'neigh_op_rgt_2')
// (4, 15, 'neigh_op_bnr_2')
// (5, 11, 'sp4_r_v_b_40')
// (5, 12, 'local_g1_5')
// (5, 12, 'lutff_0/in_0')
// (5, 12, 'sp4_r_v_b_29')
// (5, 13, 'neigh_op_top_2')
// (5, 13, 'sp4_r_v_b_16')
// (5, 14, 'lutff_2/out')
// (5, 14, 'sp4_r_v_b_5')
// (5, 15, 'neigh_op_bot_2')
// (6, 10, 'sp4_v_t_40')
// (6, 11, 'sp4_v_b_40')
// (6, 12, 'sp4_v_b_29')
// (6, 13, 'neigh_op_tnl_2')
// (6, 13, 'sp4_v_b_16')
// (6, 14, 'neigh_op_lft_2')
// (6, 14, 'sp4_v_b_5')
// (6, 15, 'neigh_op_bnl_2')

reg n236 = 0;
// (4, 13, 'neigh_op_tnr_3')
// (4, 14, 'neigh_op_rgt_3')
// (4, 15, 'neigh_op_bnr_3')
// (5, 13, 'neigh_op_top_3')
// (5, 14, 'local_g1_3')
// (5, 14, 'lutff_2/in_0')
// (5, 14, 'lutff_3/out')
// (5, 15, 'neigh_op_bot_3')
// (6, 13, 'neigh_op_tnl_3')
// (6, 14, 'neigh_op_lft_3')
// (6, 15, 'neigh_op_bnl_3')

reg n237 = 0;
// (4, 13, 'neigh_op_tnr_5')
// (4, 14, 'neigh_op_rgt_5')
// (4, 15, 'neigh_op_bnr_5')
// (5, 13, 'neigh_op_top_5')
// (5, 14, 'local_g1_5')
// (5, 14, 'lutff_5/out')
// (5, 14, 'lutff_6/in_0')
// (5, 15, 'neigh_op_bot_5')
// (6, 13, 'neigh_op_tnl_5')
// (6, 14, 'neigh_op_lft_5')
// (6, 15, 'neigh_op_bnl_5')

reg n238 = 0;
// (4, 13, 'neigh_op_tnr_6')
// (4, 14, 'neigh_op_rgt_6')
// (4, 15, 'neigh_op_bnr_6')
// (5, 13, 'neigh_op_top_6')
// (5, 14, 'local_g1_6')
// (5, 14, 'lutff_3/in_0')
// (5, 14, 'lutff_6/out')
// (5, 15, 'neigh_op_bot_6')
// (6, 13, 'neigh_op_tnl_6')
// (6, 14, 'neigh_op_lft_6')
// (6, 15, 'neigh_op_bnl_6')

wire n239;
// (5, 0, 'logic_op_tnr_1')
// (5, 1, 'neigh_op_rgt_1')
// (5, 1, 'sp4_r_v_b_34')
// (5, 2, 'neigh_op_bnr_1')
// (5, 2, 'sp4_r_v_b_23')
// (5, 3, 'sp4_r_v_b_10')
// (6, 0, 'logic_op_top_1')
// (6, 0, 'span4_vert_34')
// (6, 1, 'lutff_1/out')
// (6, 1, 'sp4_v_b_34')
// (6, 2, 'local_g0_1')
// (6, 2, 'local_g1_1')
// (6, 2, 'lutff_0/in_2')
// (6, 2, 'lutff_7/in_2')
// (6, 2, 'neigh_op_bot_1')
// (6, 2, 'sp4_v_b_23')
// (6, 3, 'local_g0_2')
// (6, 3, 'local_g1_2')
// (6, 3, 'lutff_3/in_2')
// (6, 3, 'lutff_6/in_2')
// (6, 3, 'sp4_v_b_10')
// (7, 0, 'logic_op_tnl_1')
// (7, 1, 'neigh_op_lft_1')
// (7, 2, 'neigh_op_bnl_1')

reg n240 = 0;
// (5, 0, 'span12_vert_8')
// (5, 1, 'sp12_v_b_8')
// (5, 2, 'sp12_v_b_7')
// (5, 3, 'sp12_v_b_4')
// (5, 4, 'local_g2_3')
// (5, 4, 'lutff_6/in_3')
// (5, 4, 'sp12_v_b_3')
// (5, 5, 'sp12_h_r_0')
// (5, 5, 'sp12_v_b_0')
// (6, 5, 'sp12_h_r_3')
// (7, 5, 'sp12_h_r_4')
// (8, 5, 'sp12_h_r_7')
// (9, 5, 'sp12_h_r_8')
// (10, 4, 'neigh_op_tnr_2')
// (10, 5, 'neigh_op_rgt_2')
// (10, 5, 'sp12_h_r_11')
// (10, 6, 'neigh_op_bnr_2')
// (11, 4, 'neigh_op_top_2')
// (11, 5, 'lutff_2/out')
// (11, 5, 'sp12_h_r_12')
// (11, 6, 'neigh_op_bot_2')
// (12, 4, 'neigh_op_tnl_2')
// (12, 5, 'neigh_op_lft_2')
// (12, 5, 'sp12_h_r_15')
// (12, 6, 'neigh_op_bnl_2')
// (13, 5, 'span12_horz_15')

wire n241;
// (5, 1, 'neigh_op_tnr_0')
// (5, 2, 'local_g2_0')
// (5, 2, 'local_g3_0')
// (5, 2, 'lutff_5/in_2')
// (5, 2, 'lutff_6/in_3')
// (5, 2, 'lutff_7/in_3')
// (5, 2, 'neigh_op_rgt_0')
// (5, 3, 'neigh_op_bnr_0')
// (6, 1, 'neigh_op_top_0')
// (6, 2, 'lutff_0/out')
// (6, 3, 'neigh_op_bot_0')
// (7, 1, 'neigh_op_tnl_0')
// (7, 2, 'neigh_op_lft_0')
// (7, 3, 'neigh_op_bnl_0')

wire n242;
// (5, 1, 'neigh_op_tnr_1')
// (5, 2, 'neigh_op_rgt_1')
// (5, 3, 'neigh_op_bnr_1')
// (6, 1, 'neigh_op_top_1')
// (6, 2, 'lutff_1/out')
// (6, 3, 'neigh_op_bot_1')
// (7, 1, 'neigh_op_tnl_1')
// (7, 2, 'neigh_op_lft_1')
// (7, 3, 'local_g2_1')
// (7, 3, 'local_g3_1')
// (7, 3, 'lutff_3/in_0')
// (7, 3, 'lutff_4/in_0')
// (7, 3, 'lutff_5/in_0')
// (7, 3, 'lutff_6/in_0')
// (7, 3, 'neigh_op_bnl_1')

wire n243;
// (5, 1, 'neigh_op_tnr_2')
// (5, 1, 'sp4_r_v_b_33')
// (5, 2, 'neigh_op_rgt_2')
// (5, 2, 'sp4_r_v_b_20')
// (5, 3, 'local_g2_1')
// (5, 3, 'lutff_2/in_1')
// (5, 3, 'neigh_op_bnr_2')
// (5, 3, 'sp4_r_v_b_9')
// (6, 0, 'span4_vert_33')
// (6, 1, 'neigh_op_top_2')
// (6, 1, 'sp4_v_b_33')
// (6, 2, 'lutff_2/out')
// (6, 2, 'sp4_v_b_20')
// (6, 3, 'neigh_op_bot_2')
// (6, 3, 'sp4_v_b_9')
// (7, 1, 'neigh_op_tnl_2')
// (7, 2, 'neigh_op_lft_2')
// (7, 3, 'local_g2_2')
// (7, 3, 'lutff_1/in_1')
// (7, 3, 'neigh_op_bnl_2')

wire n244;
// (5, 1, 'neigh_op_tnr_3')
// (5, 2, 'neigh_op_rgt_3')
// (5, 3, 'neigh_op_bnr_3')
// (6, 1, 'neigh_op_top_3')
// (6, 2, 'local_g0_3')
// (6, 2, 'local_g1_3')
// (6, 2, 'lutff_0/in_0')
// (6, 2, 'lutff_3/out')
// (6, 2, 'lutff_7/in_0')
// (6, 3, 'neigh_op_bot_3')
// (7, 1, 'neigh_op_tnl_3')
// (7, 2, 'neigh_op_lft_3')
// (7, 3, 'neigh_op_bnl_3')

wire n245;
// (5, 1, 'neigh_op_tnr_4')
// (5, 2, 'neigh_op_rgt_4')
// (5, 3, 'neigh_op_bnr_4')
// (6, 1, 'neigh_op_top_4')
// (6, 2, 'local_g0_4')
// (6, 2, 'lutff_4/out')
// (6, 2, 'lutff_5/in_1')
// (6, 3, 'neigh_op_bot_4')
// (7, 1, 'neigh_op_tnl_4')
// (7, 2, 'local_g1_4')
// (7, 2, 'lutff_3/in_0')
// (7, 2, 'neigh_op_lft_4')
// (7, 3, 'neigh_op_bnl_4')

wire n246;
// (5, 1, 'neigh_op_tnr_5')
// (5, 2, 'local_g2_5')
// (5, 2, 'local_g3_5')
// (5, 2, 'lutff_5/in_1')
// (5, 2, 'lutff_7/in_2')
// (5, 2, 'neigh_op_rgt_5')
// (5, 3, 'neigh_op_bnr_5')
// (6, 1, 'neigh_op_top_5')
// (6, 2, 'local_g1_5')
// (6, 2, 'lutff_2/in_0')
// (6, 2, 'lutff_5/out')
// (6, 3, 'neigh_op_bot_5')
// (7, 1, 'neigh_op_tnl_5')
// (7, 2, 'neigh_op_lft_5')
// (7, 3, 'neigh_op_bnl_5')

wire n247;
// (5, 1, 'neigh_op_tnr_6')
// (5, 1, 'sp4_r_v_b_25')
// (5, 2, 'neigh_op_rgt_6')
// (5, 2, 'sp4_r_v_b_12')
// (5, 3, 'neigh_op_bnr_6')
// (5, 3, 'sp4_r_v_b_1')
// (6, 0, 'span4_vert_25')
// (6, 1, 'neigh_op_top_6')
// (6, 1, 'sp4_v_b_25')
// (6, 2, 'lutff_6/out')
// (6, 2, 'sp4_v_b_12')
// (6, 3, 'local_g0_1')
// (6, 3, 'local_g0_6')
// (6, 3, 'lutff_3/in_0')
// (6, 3, 'lutff_6/in_0')
// (6, 3, 'neigh_op_bot_6')
// (6, 3, 'sp4_v_b_1')
// (7, 1, 'neigh_op_tnl_6')
// (7, 2, 'neigh_op_lft_6')
// (7, 3, 'neigh_op_bnl_6')

wire n248;
// (5, 1, 'neigh_op_tnr_7')
// (5, 2, 'neigh_op_rgt_7')
// (5, 3, 'neigh_op_bnr_7')
// (6, 1, 'neigh_op_top_7')
// (6, 2, 'local_g2_7')
// (6, 2, 'lutff_2/in_3')
// (6, 2, 'lutff_7/out')
// (6, 3, 'neigh_op_bot_7')
// (7, 1, 'neigh_op_tnl_7')
// (7, 2, 'neigh_op_lft_7')
// (7, 3, 'neigh_op_bnl_7')

wire n249;
// (5, 1, 'sp4_r_v_b_31')
// (5, 2, 'sp4_r_v_b_18')
// (5, 3, 'sp4_r_v_b_7')
// (6, 0, 'span4_vert_31')
// (6, 1, 'sp4_v_b_31')
// (6, 2, 'local_g0_2')
// (6, 2, 'lutff_7/in_1')
// (6, 2, 'sp4_v_b_18')
// (6, 3, 'local_g1_7')
// (6, 3, 'lutff_3/in_3')
// (6, 3, 'sp4_h_r_2')
// (6, 3, 'sp4_v_b_7')
// (7, 2, 'neigh_op_tnr_5')
// (7, 3, 'neigh_op_rgt_5')
// (7, 3, 'sp4_h_r_15')
// (7, 4, 'neigh_op_bnr_5')
// (8, 2, 'neigh_op_top_5')
// (8, 3, 'local_g0_5')
// (8, 3, 'lutff_1/in_2')
// (8, 3, 'lutff_5/out')
// (8, 3, 'sp4_h_r_26')
// (8, 4, 'neigh_op_bot_5')
// (9, 2, 'neigh_op_tnl_5')
// (9, 3, 'neigh_op_lft_5')
// (9, 3, 'sp4_h_r_39')
// (9, 4, 'neigh_op_bnl_5')
// (10, 3, 'sp4_h_l_39')

wire n250;
// (5, 2, 'neigh_op_tnr_0')
// (5, 3, 'neigh_op_rgt_0')
// (5, 4, 'neigh_op_bnr_0')
// (6, 1, 'sp4_r_v_b_41')
// (6, 2, 'neigh_op_top_0')
// (6, 2, 'sp4_r_v_b_28')
// (6, 3, 'lutff_0/out')
// (6, 3, 'sp4_h_r_0')
// (6, 3, 'sp4_r_v_b_17')
// (6, 4, 'neigh_op_bot_0')
// (6, 4, 'sp4_r_v_b_4')
// (7, 0, 'span4_vert_41')
// (7, 1, 'sp4_v_b_41')
// (7, 2, 'neigh_op_tnl_0')
// (7, 2, 'sp4_v_b_28')
// (7, 3, 'neigh_op_lft_0')
// (7, 3, 'sp4_h_r_13')
// (7, 3, 'sp4_v_b_17')
// (7, 4, 'neigh_op_bnl_0')
// (7, 4, 'sp4_h_r_4')
// (7, 4, 'sp4_v_b_4')
// (8, 3, 'sp4_h_r_24')
// (8, 4, 'sp4_h_r_17')
// (9, 3, 'sp4_h_r_37')
// (9, 4, 'sp4_h_r_28')
// (9, 4, 'sp4_r_v_b_37')
// (9, 5, 'sp4_r_v_b_24')
// (9, 6, 'sp4_r_v_b_13')
// (9, 7, 'sp4_r_v_b_0')
// (9, 8, 'sp4_r_v_b_37')
// (9, 9, 'local_g0_0')
// (9, 9, 'lutff_7/in_1')
// (9, 9, 'sp4_r_v_b_24')
// (9, 10, 'sp4_r_v_b_13')
// (9, 11, 'sp4_r_v_b_0')
// (10, 3, 'sp4_h_l_37')
// (10, 3, 'sp4_v_t_37')
// (10, 4, 'sp4_h_r_41')
// (10, 4, 'sp4_v_b_37')
// (10, 5, 'sp4_r_v_b_44')
// (10, 5, 'sp4_v_b_24')
// (10, 6, 'sp4_r_v_b_33')
// (10, 6, 'sp4_v_b_13')
// (10, 7, 'sp4_r_v_b_20')
// (10, 7, 'sp4_v_b_0')
// (10, 7, 'sp4_v_t_37')
// (10, 8, 'sp4_r_v_b_9')
// (10, 8, 'sp4_v_b_37')
// (10, 9, 'sp4_r_v_b_37')
// (10, 9, 'sp4_v_b_24')
// (10, 10, 'sp4_r_v_b_24')
// (10, 10, 'sp4_v_b_13')
// (10, 11, 'sp4_r_v_b_13')
// (10, 11, 'sp4_v_b_0')
// (10, 12, 'sp4_r_v_b_0')
// (11, 4, 'sp4_h_l_41')
// (11, 4, 'sp4_v_t_44')
// (11, 5, 'sp4_v_b_44')
// (11, 6, 'sp4_v_b_33')
// (11, 7, 'sp4_v_b_20')
// (11, 8, 'local_g0_1')
// (11, 8, 'lutff_7/in_2')
// (11, 8, 'sp4_v_b_9')
// (11, 8, 'sp4_v_t_37')
// (11, 9, 'local_g2_5')
// (11, 9, 'lutff_4/in_1')
// (11, 9, 'sp4_v_b_37')
// (11, 10, 'sp4_v_b_24')
// (11, 11, 'sp4_v_b_13')
// (11, 12, 'sp4_v_b_0')

wire n251;
// (5, 2, 'neigh_op_tnr_1')
// (5, 3, 'neigh_op_rgt_1')
// (5, 4, 'neigh_op_bnr_1')
// (6, 2, 'neigh_op_top_1')
// (6, 3, 'local_g1_1')
// (6, 3, 'lutff_1/out')
// (6, 3, 'lutff_4/in_2')
// (6, 4, 'neigh_op_bot_1')
// (7, 2, 'neigh_op_tnl_1')
// (7, 3, 'local_g0_1')
// (7, 3, 'lutff_0/in_1')
// (7, 3, 'neigh_op_lft_1')
// (7, 4, 'neigh_op_bnl_1')

wire n252;
// (5, 2, 'neigh_op_tnr_2')
// (5, 3, 'local_g3_2')
// (5, 3, 'lutff_4/in_1')
// (5, 3, 'neigh_op_rgt_2')
// (5, 4, 'neigh_op_bnr_2')
// (6, 2, 'neigh_op_top_2')
// (6, 3, 'lutff_2/out')
// (6, 4, 'neigh_op_bot_2')
// (7, 2, 'neigh_op_tnl_2')
// (7, 3, 'neigh_op_lft_2')
// (7, 4, 'neigh_op_bnl_2')

wire n253;
// (5, 2, 'neigh_op_tnr_3')
// (5, 3, 'neigh_op_rgt_3')
// (5, 4, 'neigh_op_bnr_3')
// (6, 2, 'neigh_op_top_3')
// (6, 3, 'local_g1_3')
// (6, 3, 'lutff_1/in_3')
// (6, 3, 'lutff_3/out')
// (6, 4, 'neigh_op_bot_3')
// (7, 2, 'neigh_op_tnl_3')
// (7, 3, 'neigh_op_lft_3')
// (7, 4, 'neigh_op_bnl_3')

wire n254;
// (5, 2, 'neigh_op_tnr_4')
// (5, 3, 'neigh_op_rgt_4')
// (5, 4, 'neigh_op_bnr_4')
// (6, 2, 'neigh_op_top_4')
// (6, 3, 'local_g0_4')
// (6, 3, 'lutff_0/in_0')
// (6, 3, 'lutff_4/out')
// (6, 4, 'neigh_op_bot_4')
// (7, 2, 'neigh_op_tnl_4')
// (7, 3, 'neigh_op_lft_4')
// (7, 4, 'neigh_op_bnl_4')

wire n255;
// (5, 2, 'neigh_op_tnr_5')
// (5, 3, 'neigh_op_rgt_5')
// (5, 4, 'neigh_op_bnr_5')
// (6, 2, 'neigh_op_top_5')
// (6, 3, 'local_g0_5')
// (6, 3, 'lutff_0/in_1')
// (6, 3, 'lutff_5/out')
// (6, 4, 'neigh_op_bot_5')
// (7, 2, 'neigh_op_tnl_5')
// (7, 3, 'neigh_op_lft_5')
// (7, 4, 'neigh_op_bnl_5')

wire n256;
// (5, 2, 'neigh_op_tnr_6')
// (5, 3, 'neigh_op_rgt_6')
// (5, 4, 'neigh_op_bnr_6')
// (6, 2, 'neigh_op_top_6')
// (6, 2, 'sp4_r_v_b_40')
// (6, 3, 'local_g1_5')
// (6, 3, 'local_g3_6')
// (6, 3, 'lutff_5/in_3')
// (6, 3, 'lutff_6/out')
// (6, 3, 'lutff_7/in_2')
// (6, 3, 'sp4_r_v_b_29')
// (6, 4, 'neigh_op_bot_6')
// (6, 4, 'sp4_r_v_b_16')
// (6, 5, 'sp4_r_v_b_5')
// (7, 1, 'sp4_v_t_40')
// (7, 2, 'neigh_op_tnl_6')
// (7, 2, 'sp4_v_b_40')
// (7, 3, 'neigh_op_lft_6')
// (7, 3, 'sp4_v_b_29')
// (7, 4, 'neigh_op_bnl_6')
// (7, 4, 'sp4_v_b_16')
// (7, 5, 'sp4_v_b_5')

wire n257;
// (5, 2, 'sp4_h_r_11')
// (5, 3, 'sp4_h_r_2')
// (6, 2, 'local_g1_6')
// (6, 2, 'lutff_0/in_3')
// (6, 2, 'sp4_h_r_22')
// (6, 3, 'local_g0_7')
// (6, 3, 'lutff_6/in_1')
// (6, 3, 'sp4_h_r_15')
// (7, 2, 'sp4_h_r_35')
// (7, 3, 'neigh_op_tnr_6')
// (7, 3, 'sp4_h_r_26')
// (7, 4, 'neigh_op_rgt_6')
// (7, 5, 'neigh_op_bnr_6')
// (8, 0, 'span12_vert_19')
// (8, 1, 'sp12_v_b_19')
// (8, 2, 'local_g2_0')
// (8, 2, 'lutff_1/in_1')
// (8, 2, 'lutff_7/in_3')
// (8, 2, 'sp12_v_b_16')
// (8, 2, 'sp4_h_r_46')
// (8, 3, 'neigh_op_top_6')
// (8, 3, 'sp12_v_b_15')
// (8, 3, 'sp4_h_r_39')
// (8, 3, 'sp4_r_v_b_40')
// (8, 4, 'lutff_6/out')
// (8, 4, 'sp12_v_b_12')
// (8, 4, 'sp4_r_v_b_29')
// (8, 4, 'sp4_r_v_b_45')
// (8, 5, 'neigh_op_bot_6')
// (8, 5, 'sp12_v_b_11')
// (8, 5, 'sp4_r_v_b_16')
// (8, 5, 'sp4_r_v_b_32')
// (8, 6, 'sp12_v_b_8')
// (8, 6, 'sp4_r_v_b_21')
// (8, 6, 'sp4_r_v_b_5')
// (8, 7, 'sp12_v_b_7')
// (8, 7, 'sp4_r_v_b_8')
// (8, 8, 'sp12_v_b_4')
// (8, 9, 'sp12_v_b_3')
// (8, 10, 'sp12_v_b_0')
// (9, 2, 'sp4_h_l_46')
// (9, 2, 'sp4_v_t_40')
// (9, 3, 'neigh_op_tnl_6')
// (9, 3, 'sp4_h_l_39')
// (9, 3, 'sp4_v_b_40')
// (9, 3, 'sp4_v_t_45')
// (9, 4, 'neigh_op_lft_6')
// (9, 4, 'sp4_v_b_29')
// (9, 4, 'sp4_v_b_45')
// (9, 5, 'neigh_op_bnl_6')
// (9, 5, 'sp4_v_b_16')
// (9, 5, 'sp4_v_b_32')
// (9, 6, 'sp4_v_b_21')
// (9, 6, 'sp4_v_b_5')
// (9, 7, 'sp4_v_b_8')

wire n258;
// (5, 3, 'neigh_op_tnr_2')
// (5, 4, 'neigh_op_rgt_2')
// (5, 4, 'sp4_r_v_b_36')
// (5, 5, 'local_g1_1')
// (5, 5, 'local_g1_2')
// (5, 5, 'lutff_2/in_0')
// (5, 5, 'lutff_3/in_0')
// (5, 5, 'neigh_op_bnr_2')
// (5, 5, 'sp4_r_v_b_25')
// (5, 6, 'sp4_r_v_b_12')
// (5, 7, 'sp4_r_v_b_1')
// (6, 3, 'neigh_op_top_2')
// (6, 3, 'sp4_v_t_36')
// (6, 4, 'lutff_2/out')
// (6, 4, 'sp4_v_b_36')
// (6, 5, 'neigh_op_bot_2')
// (6, 5, 'sp4_v_b_25')
// (6, 6, 'sp4_v_b_12')
// (6, 7, 'sp4_v_b_1')
// (7, 3, 'neigh_op_tnl_2')
// (7, 4, 'neigh_op_lft_2')
// (7, 5, 'neigh_op_bnl_2')

wire n259;
// (5, 3, 'neigh_op_tnr_3')
// (5, 4, 'neigh_op_rgt_3')
// (5, 4, 'sp4_r_v_b_38')
// (5, 5, 'neigh_op_bnr_3')
// (5, 5, 'sp4_r_v_b_27')
// (5, 6, 'local_g2_6')
// (5, 6, 'lutff_4/in_0')
// (5, 6, 'lutff_7/in_1')
// (5, 6, 'sp4_r_v_b_14')
// (5, 7, 'sp4_r_v_b_3')
// (6, 3, 'neigh_op_top_3')
// (6, 3, 'sp4_v_t_38')
// (6, 4, 'lutff_3/out')
// (6, 4, 'sp4_v_b_38')
// (6, 5, 'neigh_op_bot_3')
// (6, 5, 'sp4_v_b_27')
// (6, 6, 'sp4_v_b_14')
// (6, 7, 'sp4_v_b_3')
// (7, 3, 'neigh_op_tnl_3')
// (7, 4, 'neigh_op_lft_3')
// (7, 5, 'neigh_op_bnl_3')

wire n260;
// (5, 3, 'neigh_op_tnr_4')
// (5, 4, 'neigh_op_rgt_4')
// (5, 5, 'neigh_op_bnr_4')
// (6, 3, 'neigh_op_top_4')
// (6, 4, 'lutff_4/out')
// (6, 5, 'neigh_op_bot_4')
// (7, 3, 'neigh_op_tnl_4')
// (7, 4, 'local_g0_4')
// (7, 4, 'lutff_0/in_2')
// (7, 4, 'neigh_op_lft_4')
// (7, 5, 'neigh_op_bnl_4')

wire n261;
// (5, 3, 'neigh_op_tnr_7')
// (5, 4, 'neigh_op_rgt_7')
// (5, 4, 'sp4_r_v_b_46')
// (5, 5, 'neigh_op_bnr_7')
// (5, 5, 'sp4_r_v_b_35')
// (5, 5, 'sp4_r_v_b_40')
// (5, 6, 'local_g1_5')
// (5, 6, 'local_g3_6')
// (5, 6, 'lutff_1/in_0')
// (5, 6, 'lutff_2/in_0')
// (5, 6, 'sp4_r_v_b_22')
// (5, 6, 'sp4_r_v_b_29')
// (5, 7, 'sp4_r_v_b_11')
// (5, 7, 'sp4_r_v_b_16')
// (5, 8, 'sp4_r_v_b_5')
// (6, 0, 'span12_vert_21')
// (6, 1, 'sp12_v_b_21')
// (6, 2, 'sp12_v_b_18')
// (6, 3, 'neigh_op_top_7')
// (6, 3, 'sp12_v_b_17')
// (6, 3, 'sp4_v_t_46')
// (6, 4, 'lutff_7/out')
// (6, 4, 'sp12_v_b_14')
// (6, 4, 'sp4_v_b_46')
// (6, 4, 'sp4_v_t_40')
// (6, 5, 'neigh_op_bot_7')
// (6, 5, 'sp12_v_b_13')
// (6, 5, 'sp4_v_b_35')
// (6, 5, 'sp4_v_b_40')
// (6, 6, 'sp12_v_b_10')
// (6, 6, 'sp4_v_b_22')
// (6, 6, 'sp4_v_b_29')
// (6, 7, 'sp12_v_b_9')
// (6, 7, 'sp4_v_b_11')
// (6, 7, 'sp4_v_b_16')
// (6, 8, 'sp12_v_b_6')
// (6, 8, 'sp4_v_b_5')
// (6, 9, 'sp12_v_b_5')
// (6, 10, 'sp12_v_b_2')
// (6, 11, 'sp12_v_b_1')
// (7, 3, 'neigh_op_tnl_7')
// (7, 4, 'neigh_op_lft_7')
// (7, 5, 'neigh_op_bnl_7')

wire n262;
// (5, 4, 'neigh_op_tnr_1')
// (5, 5, 'local_g3_1')
// (5, 5, 'lutff_5/in_1')
// (5, 5, 'neigh_op_rgt_1')
// (5, 6, 'local_g0_1')
// (5, 6, 'lutff_0/in_1')
// (5, 6, 'lutff_5/in_2')
// (5, 6, 'neigh_op_bnr_1')
// (6, 4, 'neigh_op_top_1')
// (6, 5, 'lutff_1/out')
// (6, 6, 'neigh_op_bot_1')
// (7, 4, 'neigh_op_tnl_1')
// (7, 5, 'neigh_op_lft_1')
// (7, 6, 'neigh_op_bnl_1')

wire n263;
// (5, 4, 'neigh_op_tnr_3')
// (5, 5, 'local_g2_3')
// (5, 5, 'local_g3_3')
// (5, 5, 'lutff_0/in_2')
// (5, 5, 'lutff_3/in_2')
// (5, 5, 'neigh_op_rgt_3')
// (5, 6, 'neigh_op_bnr_3')
// (6, 4, 'neigh_op_top_3')
// (6, 5, 'lutff_3/out')
// (6, 6, 'neigh_op_bot_3')
// (7, 4, 'neigh_op_tnl_3')
// (7, 5, 'neigh_op_lft_3')
// (7, 6, 'neigh_op_bnl_3')

wire n264;
// (5, 4, 'neigh_op_tnr_4')
// (5, 5, 'neigh_op_rgt_4')
// (5, 6, 'neigh_op_bnr_4')
// (6, 4, 'neigh_op_top_4')
// (6, 5, 'local_g0_4')
// (6, 5, 'local_g1_4')
// (6, 5, 'lutff_0/in_1')
// (6, 5, 'lutff_1/in_1')
// (6, 5, 'lutff_2/in_1')
// (6, 5, 'lutff_3/in_1')
// (6, 5, 'lutff_4/out')
// (6, 6, 'neigh_op_bot_4')
// (7, 4, 'neigh_op_tnl_4')
// (7, 5, 'neigh_op_lft_4')
// (7, 6, 'neigh_op_bnl_4')

wire n265;
// (5, 4, 'neigh_op_tnr_5')
// (5, 5, 'local_g2_5')
// (5, 5, 'local_g3_5')
// (5, 5, 'lutff_1/in_2')
// (5, 5, 'lutff_2/in_2')
// (5, 5, 'lutff_4/in_2')
// (5, 5, 'lutff_6/in_3')
// (5, 5, 'neigh_op_rgt_5')
// (5, 6, 'neigh_op_bnr_5')
// (6, 4, 'neigh_op_top_5')
// (6, 5, 'lutff_5/out')
// (6, 6, 'neigh_op_bot_5')
// (7, 4, 'neigh_op_tnl_5')
// (7, 5, 'neigh_op_lft_5')
// (7, 6, 'neigh_op_bnl_5')

wire n266;
// (5, 4, 'neigh_op_tnr_6')
// (5, 5, 'local_g2_6')
// (5, 5, 'local_g3_6')
// (5, 5, 'lutff_1/in_0')
// (5, 5, 'lutff_4/in_0')
// (5, 5, 'neigh_op_rgt_6')
// (5, 6, 'neigh_op_bnr_6')
// (6, 4, 'neigh_op_top_6')
// (6, 5, 'lutff_6/out')
// (6, 6, 'neigh_op_bot_6')
// (7, 4, 'neigh_op_tnl_6')
// (7, 5, 'neigh_op_lft_6')
// (7, 6, 'neigh_op_bnl_6')

wire n267;
// (5, 4, 'neigh_op_tnr_7')
// (5, 5, 'neigh_op_rgt_7')
// (5, 6, 'neigh_op_bnr_7')
// (6, 4, 'neigh_op_top_7')
// (6, 5, 'local_g0_7')
// (6, 5, 'local_g1_7')
// (6, 5, 'lutff_0/in_0')
// (6, 5, 'lutff_1/in_0')
// (6, 5, 'lutff_2/in_0')
// (6, 5, 'lutff_3/in_0')
// (6, 5, 'lutff_7/out')
// (6, 6, 'neigh_op_bot_7')
// (7, 4, 'neigh_op_tnl_7')
// (7, 5, 'neigh_op_lft_7')
// (7, 6, 'neigh_op_bnl_7')

wire n268;
// (5, 4, 'sp4_h_r_8')
// (6, 3, 'neigh_op_tnr_0')
// (6, 4, 'neigh_op_rgt_0')
// (6, 4, 'sp4_h_r_21')
// (6, 5, 'neigh_op_bnr_0')
// (7, 0, 'span12_vert_23')
// (7, 1, 'sp12_v_b_23')
// (7, 2, 'sp12_v_b_20')
// (7, 3, 'neigh_op_top_0')
// (7, 3, 'sp12_v_b_19')
// (7, 4, 'lutff_0/out')
// (7, 4, 'sp12_v_b_16')
// (7, 4, 'sp4_h_r_32')
// (7, 5, 'neigh_op_bot_0')
// (7, 5, 'sp12_v_b_15')
// (7, 6, 'local_g3_4')
// (7, 6, 'lutff_7/in_0')
// (7, 6, 'sp12_v_b_12')
// (7, 7, 'sp12_v_b_11')
// (7, 8, 'sp12_v_b_8')
// (7, 9, 'sp12_v_b_7')
// (7, 10, 'sp12_v_b_4')
// (7, 11, 'sp12_v_b_3')
// (7, 12, 'sp12_v_b_0')
// (8, 3, 'neigh_op_tnl_0')
// (8, 4, 'neigh_op_lft_0')
// (8, 4, 'sp4_h_r_45')
// (8, 5, 'neigh_op_bnl_0')
// (8, 5, 'sp4_r_v_b_36')
// (8, 6, 'sp4_r_v_b_25')
// (8, 7, 'sp4_r_v_b_12')
// (8, 8, 'sp4_r_v_b_1')
// (8, 9, 'sp4_r_v_b_41')
// (8, 10, 'sp4_r_v_b_28')
// (8, 11, 'sp4_r_v_b_17')
// (8, 12, 'sp4_r_v_b_4')
// (9, 4, 'sp4_h_l_45')
// (9, 4, 'sp4_v_t_36')
// (9, 5, 'sp4_v_b_36')
// (9, 6, 'sp4_v_b_25')
// (9, 7, 'sp4_v_b_12')
// (9, 8, 'local_g0_1')
// (9, 8, 'lutff_3/in_2')
// (9, 8, 'sp4_v_b_1')
// (9, 8, 'sp4_v_t_41')
// (9, 9, 'local_g2_1')
// (9, 9, 'lutff_1/in_2')
// (9, 9, 'sp4_v_b_41')
// (9, 10, 'sp4_v_b_28')
// (9, 11, 'sp4_v_b_17')
// (9, 12, 'sp4_v_b_4')

wire n269;
// (5, 5, 'neigh_op_tnr_0')
// (5, 6, 'neigh_op_rgt_0')
// (5, 7, 'neigh_op_bnr_0')
// (6, 5, 'local_g0_0')
// (6, 5, 'local_g1_0')
// (6, 5, 'lutff_0/in_2')
// (6, 5, 'lutff_3/in_2')
// (6, 5, 'neigh_op_top_0')
// (6, 6, 'lutff_0/out')
// (6, 7, 'neigh_op_bot_0')
// (7, 5, 'local_g2_0')
// (7, 5, 'local_g3_0')
// (7, 5, 'lutff_1/in_0')
// (7, 5, 'lutff_5/in_0')
// (7, 5, 'lutff_6/in_2')
// (7, 5, 'neigh_op_tnl_0')
// (7, 6, 'neigh_op_lft_0')
// (7, 7, 'neigh_op_bnl_0')

wire n270;
// (5, 5, 'neigh_op_tnr_1')
// (5, 6, 'neigh_op_rgt_1')
// (5, 7, 'neigh_op_bnr_1')
// (6, 5, 'local_g0_1')
// (6, 5, 'local_g1_1')
// (6, 5, 'lutff_1/in_2')
// (6, 5, 'lutff_2/in_2')
// (6, 5, 'neigh_op_top_1')
// (6, 6, 'lutff_1/out')
// (6, 7, 'neigh_op_bot_1')
// (7, 5, 'local_g2_1')
// (7, 5, 'local_g3_1')
// (7, 5, 'lutff_1/in_1')
// (7, 5, 'lutff_5/in_1')
// (7, 5, 'lutff_6/in_3')
// (7, 5, 'neigh_op_tnl_1')
// (7, 6, 'neigh_op_lft_1')
// (7, 7, 'neigh_op_bnl_1')

wire n271;
// (5, 5, 'neigh_op_tnr_2')
// (5, 6, 'local_g1_1')
// (5, 6, 'local_g3_2')
// (5, 6, 'lutff_2/in_1')
// (5, 6, 'lutff_7/in_3')
// (5, 6, 'neigh_op_rgt_2')
// (5, 6, 'sp4_h_r_9')
// (5, 7, 'neigh_op_bnr_2')
// (6, 5, 'neigh_op_top_2')
// (6, 6, 'lutff_2/out')
// (6, 6, 'sp4_h_r_20')
// (6, 7, 'neigh_op_bot_2')
// (7, 5, 'neigh_op_tnl_2')
// (7, 6, 'local_g0_2')
// (7, 6, 'local_g2_1')
// (7, 6, 'lutff_1/in_3')
// (7, 6, 'lutff_3/in_0')
// (7, 6, 'lutff_6/in_0')
// (7, 6, 'neigh_op_lft_2')
// (7, 6, 'sp4_h_r_33')
// (7, 7, 'neigh_op_bnl_2')
// (8, 6, 'sp4_h_r_44')
// (9, 6, 'sp4_h_l_44')

wire n272;
// (5, 5, 'neigh_op_tnr_4')
// (5, 6, 'local_g3_4')
// (5, 6, 'lutff_2/in_3')
// (5, 6, 'lutff_7/in_0')
// (5, 6, 'neigh_op_rgt_4')
// (5, 7, 'neigh_op_bnr_4')
// (6, 5, 'neigh_op_top_4')
// (6, 6, 'local_g0_4')
// (6, 6, 'lutff_4/out')
// (6, 6, 'lutff_6/in_0')
// (6, 7, 'neigh_op_bot_4')
// (7, 5, 'neigh_op_tnl_4')
// (7, 6, 'local_g0_4')
// (7, 6, 'lutff_1/in_1')
// (7, 6, 'lutff_3/in_3')
// (7, 6, 'neigh_op_lft_4')
// (7, 7, 'neigh_op_bnl_4')

wire n273;
// (5, 5, 'neigh_op_tnr_5')
// (5, 6, 'neigh_op_rgt_5')
// (5, 7, 'neigh_op_bnr_5')
// (6, 3, 'sp4_r_v_b_46')
// (6, 4, 'sp4_r_v_b_35')
// (6, 5, 'neigh_op_top_5')
// (6, 5, 'sp4_r_v_b_22')
// (6, 6, 'local_g1_5')
// (6, 6, 'lutff_1/in_1')
// (6, 6, 'lutff_2/in_2')
// (6, 6, 'lutff_5/out')
// (6, 6, 'sp4_r_v_b_11')
// (6, 7, 'neigh_op_bot_5')
// (7, 2, 'sp4_v_t_46')
// (7, 3, 'sp4_v_b_46')
// (7, 4, 'sp4_v_b_35')
// (7, 5, 'neigh_op_tnl_5')
// (7, 5, 'sp4_v_b_22')
// (7, 6, 'local_g0_3')
// (7, 6, 'local_g1_5')
// (7, 6, 'lutff_4/in_3')
// (7, 6, 'lutff_5/in_3')
// (7, 6, 'neigh_op_lft_5')
// (7, 6, 'sp4_v_b_11')
// (7, 7, 'neigh_op_bnl_5')

wire n274;
// (5, 5, 'neigh_op_tnr_6')
// (5, 6, 'neigh_op_rgt_6')
// (5, 7, 'neigh_op_bnr_6')
// (6, 5, 'local_g0_6')
// (6, 5, 'local_g1_6')
// (6, 5, 'lutff_1/in_3')
// (6, 5, 'lutff_2/in_3')
// (6, 5, 'neigh_op_top_6')
// (6, 6, 'lutff_6/out')
// (6, 7, 'neigh_op_bot_6')
// (7, 5, 'local_g3_6')
// (7, 5, 'lutff_0/in_1')
// (7, 5, 'lutff_3/in_0')
// (7, 5, 'lutff_5/in_2')
// (7, 5, 'neigh_op_tnl_6')
// (7, 6, 'neigh_op_lft_6')
// (7, 7, 'neigh_op_bnl_6')

wire n275;
// (5, 5, 'neigh_op_tnr_7')
// (5, 6, 'local_g2_7')
// (5, 6, 'local_g3_7')
// (5, 6, 'lutff_1/in_3')
// (5, 6, 'lutff_4/in_1')
// (5, 6, 'neigh_op_rgt_7')
// (5, 7, 'neigh_op_bnr_7')
// (6, 5, 'neigh_op_top_7')
// (6, 6, 'lutff_7/out')
// (6, 7, 'neigh_op_bot_7')
// (7, 5, 'neigh_op_tnl_7')
// (7, 6, 'local_g0_7')
// (7, 6, 'lutff_1/in_2')
// (7, 6, 'lutff_4/in_1')
// (7, 6, 'neigh_op_lft_7')
// (7, 7, 'neigh_op_bnl_7')

wire n276;
// (5, 6, 'neigh_op_tnr_0')
// (5, 7, 'neigh_op_rgt_0')
// (5, 8, 'neigh_op_bnr_0')
// (6, 6, 'local_g1_0')
// (6, 6, 'lutff_1/in_2')
// (6, 6, 'lutff_2/in_3')
// (6, 6, 'neigh_op_top_0')
// (6, 7, 'lutff_0/out')
// (6, 8, 'neigh_op_bot_0')
// (7, 6, 'neigh_op_tnl_0')
// (7, 7, 'neigh_op_lft_0')
// (7, 8, 'neigh_op_bnl_0')

wire n277;
// (5, 6, 'neigh_op_tnr_1')
// (5, 7, 'neigh_op_rgt_1')
// (5, 8, 'neigh_op_bnr_1')
// (6, 6, 'neigh_op_top_1')
// (6, 7, 'local_g2_1')
// (6, 7, 'lutff_1/out')
// (6, 7, 'lutff_4/in_3')
// (6, 8, 'neigh_op_bot_1')
// (7, 6, 'neigh_op_tnl_1')
// (7, 7, 'neigh_op_lft_1')
// (7, 8, 'neigh_op_bnl_1')

wire n278;
// (5, 6, 'neigh_op_tnr_2')
// (5, 7, 'neigh_op_rgt_2')
// (5, 8, 'neigh_op_bnr_2')
// (6, 6, 'local_g0_2')
// (6, 6, 'lutff_4/in_2')
// (6, 6, 'lutff_5/in_1')
// (6, 6, 'lutff_7/in_1')
// (6, 6, 'neigh_op_top_2')
// (6, 7, 'lutff_2/out')
// (6, 8, 'neigh_op_bot_2')
// (7, 6, 'local_g3_2')
// (7, 6, 'lutff_0/in_1')
// (7, 6, 'lutff_2/in_1')
// (7, 6, 'neigh_op_tnl_2')
// (7, 7, 'neigh_op_lft_2')
// (7, 8, 'neigh_op_bnl_2')

wire n279;
// (5, 6, 'neigh_op_tnr_3')
// (5, 7, 'neigh_op_rgt_3')
// (5, 8, 'neigh_op_bnr_3')
// (6, 6, 'local_g0_3')
// (6, 6, 'local_g1_3')
// (6, 6, 'lutff_3/in_3')
// (6, 6, 'lutff_6/in_3')
// (6, 6, 'neigh_op_top_3')
// (6, 7, 'lutff_3/out')
// (6, 8, 'neigh_op_bot_3')
// (7, 6, 'neigh_op_tnl_3')
// (7, 7, 'neigh_op_lft_3')
// (7, 8, 'neigh_op_bnl_3')

wire n280;
// (5, 6, 'neigh_op_tnr_4')
// (5, 7, 'neigh_op_rgt_4')
// (5, 8, 'neigh_op_bnr_4')
// (6, 6, 'neigh_op_top_4')
// (6, 7, 'local_g3_4')
// (6, 7, 'lutff_2/in_3')
// (6, 7, 'lutff_4/out')
// (6, 8, 'neigh_op_bot_4')
// (7, 6, 'neigh_op_tnl_4')
// (7, 7, 'neigh_op_lft_4')
// (7, 8, 'neigh_op_bnl_4')

reg n281 = 0;
// (5, 6, 'neigh_op_tnr_5')
// (5, 7, 'local_g2_5')
// (5, 7, 'lutff_3/in_0')
// (5, 7, 'neigh_op_rgt_5')
// (5, 8, 'neigh_op_bnr_5')
// (6, 6, 'neigh_op_top_5')
// (6, 7, 'lutff_5/out')
// (6, 8, 'neigh_op_bot_5')
// (7, 6, 'neigh_op_tnl_5')
// (7, 7, 'neigh_op_lft_5')
// (7, 8, 'neigh_op_bnl_5')

reg n282 = 0;
// (5, 6, 'neigh_op_tnr_7')
// (5, 7, 'neigh_op_rgt_7')
// (5, 8, 'neigh_op_bnr_7')
// (6, 6, 'neigh_op_top_7')
// (6, 7, 'local_g0_7')
// (6, 7, 'lutff_5/in_0')
// (6, 7, 'lutff_7/out')
// (6, 8, 'neigh_op_bot_7')
// (7, 6, 'neigh_op_tnl_7')
// (7, 7, 'neigh_op_lft_7')
// (7, 8, 'neigh_op_bnl_7')

reg n283 = 0;
// (5, 6, 'sp4_h_r_6')
// (5, 7, 'sp4_h_r_11')
// (6, 6, 'sp4_h_r_19')
// (6, 7, 'sp4_h_r_22')
// (7, 5, 'sp4_r_v_b_44')
// (7, 6, 'sp4_h_r_30')
// (7, 6, 'sp4_r_v_b_33')
// (7, 7, 'sp4_h_r_35')
// (7, 7, 'sp4_r_v_b_20')
// (7, 8, 'sp4_r_v_b_9')
// (8, 3, 'neigh_op_tnr_7')
// (8, 3, 'sp4_r_v_b_43')
// (8, 4, 'neigh_op_rgt_7')
// (8, 4, 'sp4_h_r_3')
// (8, 4, 'sp4_r_v_b_30')
// (8, 4, 'sp4_r_v_b_46')
// (8, 4, 'sp4_v_t_44')
// (8, 5, 'local_g3_3')
// (8, 5, 'local_g3_4')
// (8, 5, 'lutff_0/in_1')
// (8, 5, 'lutff_1/in_1')
// (8, 5, 'lutff_3/in_1')
// (8, 5, 'neigh_op_bnr_7')
// (8, 5, 'sp4_r_v_b_19')
// (8, 5, 'sp4_r_v_b_35')
// (8, 5, 'sp4_v_b_44')
// (8, 6, 'local_g3_3')
// (8, 6, 'local_g3_6')
// (8, 6, 'lutff_0/in_1')
// (8, 6, 'lutff_1/in_1')
// (8, 6, 'lutff_2/in_1')
// (8, 6, 'lutff_3/in_1')
// (8, 6, 'lutff_4/in_1')
// (8, 6, 'sp4_h_r_43')
// (8, 6, 'sp4_r_v_b_22')
// (8, 6, 'sp4_r_v_b_6')
// (8, 6, 'sp4_v_b_33')
// (8, 7, 'local_g2_3')
// (8, 7, 'local_g2_6')
// (8, 7, 'lutff_0/in_2')
// (8, 7, 'lutff_1/in_1')
// (8, 7, 'lutff_3/in_1')
// (8, 7, 'lutff_4/in_1')
// (8, 7, 'sp4_h_r_46')
// (8, 7, 'sp4_r_v_b_11')
// (8, 7, 'sp4_v_b_20')
// (8, 8, 'sp4_v_b_9')
// (9, 2, 'sp4_v_t_43')
// (9, 3, 'neigh_op_top_7')
// (9, 3, 'sp4_v_b_43')
// (9, 3, 'sp4_v_t_46')
// (9, 4, 'local_g0_7')
// (9, 4, 'local_g1_7')
// (9, 4, 'lutff_1/in_1')
// (9, 4, 'lutff_5/in_2')
// (9, 4, 'lutff_7/out')
// (9, 4, 'sp4_h_r_14')
// (9, 4, 'sp4_v_b_30')
// (9, 4, 'sp4_v_b_46')
// (9, 5, 'neigh_op_bot_7')
// (9, 5, 'sp4_v_b_19')
// (9, 5, 'sp4_v_b_35')
// (9, 6, 'sp4_h_l_43')
// (9, 6, 'sp4_v_b_22')
// (9, 6, 'sp4_v_b_6')
// (9, 7, 'sp4_h_l_46')
// (9, 7, 'sp4_v_b_11')
// (10, 3, 'neigh_op_tnl_7')
// (10, 4, 'neigh_op_lft_7')
// (10, 4, 'sp4_h_r_27')
// (10, 5, 'neigh_op_bnl_7')
// (11, 4, 'local_g3_6')
// (11, 4, 'lutff_6/in_1')
// (11, 4, 'sp4_h_r_38')
// (11, 5, 'sp4_r_v_b_38')
// (11, 6, 'local_g0_3')
// (11, 6, 'lutff_2/in_1')
// (11, 6, 'lutff_4/in_1')
// (11, 6, 'sp4_r_v_b_27')
// (11, 7, 'sp4_r_v_b_14')
// (11, 8, 'sp4_r_v_b_3')
// (12, 4, 'sp4_h_l_38')
// (12, 4, 'sp4_v_t_38')
// (12, 5, 'sp4_v_b_38')
// (12, 6, 'sp4_v_b_27')
// (12, 7, 'sp4_v_b_14')
// (12, 8, 'sp4_v_b_3')

wire n284;
// (5, 6, 'sp4_r_v_b_37')
// (5, 7, 'sp4_r_v_b_24')
// (5, 8, 'neigh_op_tnr_0')
// (5, 8, 'sp4_r_v_b_13')
// (5, 9, 'neigh_op_rgt_0')
// (5, 9, 'sp4_r_v_b_0')
// (5, 10, 'neigh_op_bnr_0')
// (6, 5, 'sp4_v_t_37')
// (6, 6, 'sp4_v_b_37')
// (6, 7, 'sp4_v_b_24')
// (6, 8, 'local_g1_5')
// (6, 8, 'lutff_1/in_3')
// (6, 8, 'neigh_op_top_0')
// (6, 8, 'sp4_v_b_13')
// (6, 9, 'lutff_0/out')
// (6, 9, 'sp4_v_b_0')
// (6, 10, 'neigh_op_bot_0')
// (7, 8, 'neigh_op_tnl_0')
// (7, 9, 'neigh_op_lft_0')
// (7, 10, 'neigh_op_bnl_0')

wire n285;
// (5, 7, 'neigh_op_tnr_1')
// (5, 8, 'neigh_op_rgt_1')
// (5, 9, 'neigh_op_bnr_1')
// (6, 7, 'neigh_op_top_1')
// (6, 8, 'local_g1_1')
// (6, 8, 'lutff_1/out')
// (6, 8, 'lutff_3/in_3')
// (6, 9, 'neigh_op_bot_1')
// (7, 7, 'neigh_op_tnl_1')
// (7, 8, 'neigh_op_lft_1')
// (7, 9, 'neigh_op_bnl_1')

wire n286;
// (5, 7, 'neigh_op_tnr_3')
// (5, 8, 'neigh_op_rgt_3')
// (5, 9, 'neigh_op_bnr_3')
// (6, 5, 'sp4_r_v_b_42')
// (6, 6, 'local_g0_7')
// (6, 6, 'lutff_4/in_1')
// (6, 6, 'lutff_7/in_0')
// (6, 6, 'sp4_r_v_b_31')
// (6, 7, 'neigh_op_top_3')
// (6, 7, 'sp4_r_v_b_18')
// (6, 8, 'lutff_3/out')
// (6, 8, 'sp4_r_v_b_7')
// (6, 9, 'neigh_op_bot_3')
// (7, 4, 'sp4_v_t_42')
// (7, 5, 'sp4_v_b_42')
// (7, 6, 'local_g3_7')
// (7, 6, 'lutff_0/in_0')
// (7, 6, 'lutff_2/in_0')
// (7, 6, 'sp4_v_b_31')
// (7, 7, 'local_g2_3')
// (7, 7, 'lutff_0/in_1')
// (7, 7, 'neigh_op_tnl_3')
// (7, 7, 'sp4_v_b_18')
// (7, 8, 'neigh_op_lft_3')
// (7, 8, 'sp4_v_b_7')
// (7, 9, 'neigh_op_bnl_3')

reg n287 = 0;
// (5, 7, 'neigh_op_tnr_4')
// (5, 8, 'neigh_op_rgt_4')
// (5, 8, 'sp4_r_v_b_40')
// (5, 9, 'neigh_op_bnr_4')
// (5, 9, 'sp4_r_v_b_29')
// (5, 10, 'sp4_r_v_b_16')
// (5, 11, 'sp4_r_v_b_5')
// (6, 7, 'neigh_op_top_4')
// (6, 7, 'sp4_v_t_40')
// (6, 8, 'lutff_4/out')
// (6, 8, 'sp4_v_b_40')
// (6, 9, 'local_g2_5')
// (6, 9, 'lutff_4/in_1')
// (6, 9, 'neigh_op_bot_4')
// (6, 9, 'sp4_v_b_29')
// (6, 10, 'sp4_v_b_16')
// (6, 11, 'sp4_v_b_5')
// (7, 7, 'neigh_op_tnl_4')
// (7, 8, 'neigh_op_lft_4')
// (7, 9, 'neigh_op_bnl_4')

reg n288 = 0;
// (5, 7, 'neigh_op_tnr_6')
// (5, 8, 'neigh_op_rgt_6')
// (5, 9, 'neigh_op_bnr_6')
// (6, 7, 'neigh_op_top_6')
// (6, 8, 'lutff_6/out')
// (6, 9, 'neigh_op_bot_6')
// (7, 7, 'neigh_op_tnl_6')
// (7, 8, 'local_g0_6')
// (7, 8, 'lutff_1/in_1')
// (7, 8, 'neigh_op_lft_6')
// (7, 9, 'neigh_op_bnl_6')

reg n289 = 0;
// (5, 7, 'neigh_op_tnr_7')
// (5, 8, 'neigh_op_rgt_7')
// (5, 9, 'neigh_op_bnr_7')
// (6, 7, 'neigh_op_top_7')
// (6, 8, 'lutff_7/out')
// (6, 8, 'sp4_r_v_b_47')
// (6, 9, 'neigh_op_bot_7')
// (6, 9, 'sp4_r_v_b_34')
// (6, 10, 'sp4_r_v_b_23')
// (6, 11, 'local_g2_2')
// (6, 11, 'lutff_3/in_1')
// (6, 11, 'sp4_r_v_b_10')
// (7, 7, 'neigh_op_tnl_7')
// (7, 7, 'sp4_v_t_47')
// (7, 8, 'neigh_op_lft_7')
// (7, 8, 'sp4_v_b_47')
// (7, 9, 'neigh_op_bnl_7')
// (7, 9, 'sp4_v_b_34')
// (7, 10, 'sp4_v_b_23')
// (7, 11, 'sp4_v_b_10')

reg n290 = 0;
// (5, 7, 'sp12_h_r_0')
// (6, 7, 'sp12_h_r_3')
// (7, 7, 'sp12_h_r_4')
// (8, 6, 'neigh_op_tnr_0')
// (8, 7, 'neigh_op_rgt_0')
// (8, 7, 'sp12_h_r_7')
// (8, 8, 'neigh_op_bnr_0')
// (9, 6, 'neigh_op_top_0')
// (9, 7, 'lutff_0/out')
// (9, 7, 'sp12_h_r_8')
// (9, 8, 'neigh_op_bot_0')
// (10, 6, 'neigh_op_tnl_0')
// (10, 7, 'neigh_op_lft_0')
// (10, 7, 'sp12_h_r_11')
// (10, 8, 'neigh_op_bnl_0')
// (11, 7, 'local_g1_4')
// (11, 7, 'lutff_3/in_0')
// (11, 7, 'sp12_h_r_12')
// (12, 7, 'sp12_h_r_15')
// (13, 7, 'span12_horz_15')

wire n291;
// (5, 7, 'sp4_h_r_3')
// (6, 7, 'local_g0_6')
// (6, 7, 'lutff_0/in_2')
// (6, 7, 'sp4_h_r_14')
// (7, 6, 'sp4_r_v_b_37')
// (7, 7, 'local_g1_0')
// (7, 7, 'lutff_0/in_3')
// (7, 7, 'sp4_h_r_27')
// (7, 7, 'sp4_r_v_b_24')
// (7, 8, 'neigh_op_tnr_0')
// (7, 8, 'sp4_r_v_b_13')
// (7, 9, 'neigh_op_rgt_0')
// (7, 9, 'sp4_r_v_b_0')
// (7, 10, 'neigh_op_bnr_0')
// (8, 5, 'sp4_v_t_37')
// (8, 6, 'sp4_v_b_37')
// (8, 7, 'sp4_h_r_38')
// (8, 7, 'sp4_v_b_24')
// (8, 8, 'neigh_op_top_0')
// (8, 8, 'sp4_r_v_b_44')
// (8, 8, 'sp4_v_b_13')
// (8, 9, 'lutff_0/out')
// (8, 9, 'sp4_r_v_b_33')
// (8, 9, 'sp4_v_b_0')
// (8, 10, 'neigh_op_bot_0')
// (8, 10, 'sp4_r_v_b_20')
// (8, 11, 'sp4_r_v_b_9')
// (9, 7, 'sp4_h_l_38')
// (9, 7, 'sp4_v_t_44')
// (9, 8, 'neigh_op_tnl_0')
// (9, 8, 'sp4_v_b_44')
// (9, 9, 'neigh_op_lft_0')
// (9, 9, 'sp4_v_b_33')
// (9, 10, 'neigh_op_bnl_0')
// (9, 10, 'sp4_v_b_20')
// (9, 11, 'sp4_v_b_9')

wire n292;
// (5, 7, 'sp4_r_v_b_37')
// (5, 8, 'sp4_r_v_b_24')
// (5, 9, 'neigh_op_tnr_0')
// (5, 9, 'sp4_r_v_b_13')
// (5, 10, 'neigh_op_rgt_0')
// (5, 10, 'sp4_r_v_b_0')
// (5, 11, 'neigh_op_bnr_0')
// (6, 6, 'sp4_v_t_37')
// (6, 7, 'local_g2_5')
// (6, 7, 'local_g3_5')
// (6, 7, 'lutff_2/in_1')
// (6, 7, 'lutff_7/in_1')
// (6, 7, 'sp4_v_b_37')
// (6, 8, 'sp4_v_b_24')
// (6, 9, 'neigh_op_top_0')
// (6, 9, 'sp4_v_b_13')
// (6, 10, 'lutff_0/out')
// (6, 10, 'sp4_v_b_0')
// (6, 11, 'neigh_op_bot_0')
// (7, 9, 'neigh_op_tnl_0')
// (7, 10, 'neigh_op_lft_0')
// (7, 11, 'neigh_op_bnl_0')

wire n293;
// (5, 7, 'sp4_r_v_b_42')
// (5, 8, 'neigh_op_tnr_1')
// (5, 8, 'sp4_r_v_b_31')
// (5, 9, 'local_g2_1')
// (5, 9, 'lutff_0/in_1')
// (5, 9, 'neigh_op_rgt_1')
// (5, 9, 'sp4_r_v_b_18')
// (5, 10, 'local_g1_7')
// (5, 10, 'lutff_3/in_1')
// (5, 10, 'neigh_op_bnr_1')
// (5, 10, 'sp4_r_v_b_7')
// (6, 6, 'sp4_v_t_42')
// (6, 7, 'sp4_v_b_42')
// (6, 8, 'neigh_op_top_1')
// (6, 8, 'sp4_v_b_31')
// (6, 9, 'lutff_1/out')
// (6, 9, 'sp4_v_b_18')
// (6, 10, 'neigh_op_bot_1')
// (6, 10, 'sp4_v_b_7')
// (7, 8, 'neigh_op_tnl_1')
// (7, 9, 'neigh_op_lft_1')
// (7, 10, 'neigh_op_bnl_1')

reg n294 = 0;
// (5, 8, 'neigh_op_tnr_2')
// (5, 9, 'neigh_op_rgt_2')
// (5, 10, 'neigh_op_bnr_2')
// (6, 8, 'neigh_op_top_2')
// (6, 9, 'local_g0_2')
// (6, 9, 'lutff_1/in_1')
// (6, 9, 'lutff_2/out')
// (6, 10, 'neigh_op_bot_2')
// (7, 8, 'neigh_op_tnl_2')
// (7, 9, 'neigh_op_lft_2')
// (7, 10, 'neigh_op_bnl_2')

reg n295 = 0;
// (5, 8, 'neigh_op_tnr_3')
// (5, 9, 'neigh_op_rgt_3')
// (5, 10, 'neigh_op_bnr_3')
// (6, 8, 'local_g1_3')
// (6, 8, 'lutff_4/in_0')
// (6, 8, 'neigh_op_top_3')
// (6, 9, 'local_g3_3')
// (6, 9, 'lutff_3/out')
// (6, 9, 'lutff_5/in_1')
// (6, 10, 'neigh_op_bot_3')
// (7, 8, 'neigh_op_tnl_3')
// (7, 9, 'neigh_op_lft_3')
// (7, 10, 'neigh_op_bnl_3')

reg n296 = 0;
// (5, 8, 'neigh_op_tnr_4')
// (5, 9, 'neigh_op_rgt_4')
// (5, 10, 'neigh_op_bnr_4')
// (6, 8, 'neigh_op_top_4')
// (6, 9, 'local_g1_4')
// (6, 9, 'lutff_2/in_1')
// (6, 9, 'lutff_4/out')
// (6, 10, 'neigh_op_bot_4')
// (7, 8, 'neigh_op_tnl_4')
// (7, 9, 'neigh_op_lft_4')
// (7, 10, 'neigh_op_bnl_4')

reg n297 = 0;
// (5, 8, 'neigh_op_tnr_5')
// (5, 9, 'neigh_op_rgt_5')
// (5, 10, 'neigh_op_bnr_5')
// (6, 8, 'neigh_op_top_5')
// (6, 9, 'local_g0_5')
// (6, 9, 'local_g1_5')
// (6, 9, 'lutff_4/in_2')
// (6, 9, 'lutff_5/out')
// (6, 9, 'lutff_6/in_1')
// (6, 10, 'neigh_op_bot_5')
// (7, 8, 'neigh_op_tnl_5')
// (7, 9, 'neigh_op_lft_5')
// (7, 10, 'neigh_op_bnl_5')

reg n298 = 0;
// (5, 8, 'neigh_op_tnr_6')
// (5, 9, 'neigh_op_rgt_6')
// (5, 10, 'neigh_op_bnr_6')
// (6, 8, 'neigh_op_top_6')
// (6, 9, 'local_g0_6')
// (6, 9, 'lutff_2/in_2')
// (6, 9, 'lutff_6/out')
// (6, 9, 'lutff_7/in_1')
// (6, 10, 'neigh_op_bot_6')
// (7, 8, 'neigh_op_tnl_6')
// (7, 9, 'neigh_op_lft_6')
// (7, 10, 'neigh_op_bnl_6')

reg n299 = 0;
// (5, 8, 'neigh_op_tnr_7')
// (5, 9, 'neigh_op_rgt_7')
// (5, 10, 'neigh_op_bnr_7')
// (6, 8, 'neigh_op_top_7')
// (6, 9, 'local_g0_7')
// (6, 9, 'local_g1_7')
// (6, 9, 'lutff_1/in_2')
// (6, 9, 'lutff_3/in_1')
// (6, 9, 'lutff_7/out')
// (6, 10, 'neigh_op_bot_7')
// (7, 8, 'neigh_op_tnl_7')
// (7, 9, 'neigh_op_lft_7')
// (7, 10, 'neigh_op_bnl_7')

reg n300 = 0;
// (5, 8, 'sp4_r_v_b_38')
// (5, 9, 'neigh_op_tnr_7')
// (5, 9, 'sp4_r_v_b_27')
// (5, 10, 'neigh_op_rgt_7')
// (5, 10, 'sp4_r_v_b_14')
// (5, 11, 'neigh_op_bnr_7')
// (5, 11, 'sp4_r_v_b_3')
// (5, 12, 'sp4_r_v_b_43')
// (5, 13, 'sp4_r_v_b_30')
// (5, 14, 'sp4_r_v_b_19')
// (5, 15, 'sp4_r_v_b_6')
// (6, 7, 'sp4_v_t_38')
// (6, 8, 'sp4_v_b_38')
// (6, 9, 'neigh_op_top_7')
// (6, 9, 'sp4_v_b_27')
// (6, 10, 'local_g1_7')
// (6, 10, 'lutff_1/in_1')
// (6, 10, 'lutff_7/out')
// (6, 10, 'sp4_v_b_14')
// (6, 11, 'neigh_op_bot_7')
// (6, 11, 'sp4_v_b_3')
// (6, 11, 'sp4_v_t_43')
// (6, 12, 'sp4_v_b_43')
// (6, 13, 'sp4_v_b_30')
// (6, 14, 'local_g0_3')
// (6, 14, 'lutff_7/in_0')
// (6, 14, 'sp4_v_b_19')
// (6, 15, 'sp4_v_b_6')
// (7, 9, 'neigh_op_tnl_7')
// (7, 10, 'neigh_op_lft_7')
// (7, 11, 'neigh_op_bnl_7')

reg n301 = 0;
// (5, 9, 'neigh_op_tnr_1')
// (5, 10, 'neigh_op_rgt_1')
// (5, 11, 'neigh_op_bnr_1')
// (6, 9, 'neigh_op_top_1')
// (6, 10, 'local_g0_1')
// (6, 10, 'local_g1_1')
// (6, 10, 'lutff_1/out')
// (6, 10, 'lutff_3/in_1')
// (6, 10, 'lutff_5/in_2')
// (6, 11, 'neigh_op_bot_1')
// (7, 9, 'neigh_op_tnl_1')
// (7, 10, 'neigh_op_lft_1')
// (7, 11, 'neigh_op_bnl_1')

reg n302 = 0;
// (5, 9, 'neigh_op_tnr_2')
// (5, 10, 'neigh_op_rgt_2')
// (5, 11, 'neigh_op_bnr_2')
// (6, 9, 'neigh_op_top_2')
// (6, 10, 'local_g2_2')
// (6, 10, 'lutff_0/in_2')
// (6, 10, 'lutff_2/out')
// (6, 10, 'lutff_7/in_1')
// (6, 11, 'neigh_op_bot_2')
// (7, 9, 'neigh_op_tnl_2')
// (7, 10, 'neigh_op_lft_2')
// (7, 11, 'neigh_op_bnl_2')

reg n303 = 0;
// (5, 9, 'neigh_op_tnr_3')
// (5, 10, 'neigh_op_rgt_3')
// (5, 11, 'neigh_op_bnr_3')
// (6, 9, 'neigh_op_top_3')
// (6, 10, 'local_g0_3')
// (6, 10, 'local_g1_3')
// (6, 10, 'lutff_2/in_1')
// (6, 10, 'lutff_3/out')
// (6, 10, 'lutff_6/in_2')
// (6, 11, 'neigh_op_bot_3')
// (7, 9, 'neigh_op_tnl_3')
// (7, 10, 'neigh_op_lft_3')
// (7, 11, 'neigh_op_bnl_3')

reg n304 = 0;
// (5, 9, 'neigh_op_tnr_4')
// (5, 10, 'neigh_op_rgt_4')
// (5, 11, 'neigh_op_bnr_4')
// (6, 7, 'sp4_r_v_b_44')
// (6, 8, 'sp4_r_v_b_33')
// (6, 9, 'neigh_op_top_4')
// (6, 9, 'sp4_r_v_b_20')
// (6, 10, 'lutff_4/out')
// (6, 10, 'sp4_r_v_b_9')
// (6, 11, 'neigh_op_bot_4')
// (6, 11, 'sp4_r_v_b_44')
// (6, 12, 'local_g2_1')
// (6, 12, 'lutff_1/in_0')
// (6, 12, 'sp4_r_v_b_33')
// (6, 13, 'sp4_r_v_b_20')
// (6, 14, 'sp4_r_v_b_9')
// (7, 6, 'sp4_v_t_44')
// (7, 7, 'sp4_v_b_44')
// (7, 8, 'sp4_v_b_33')
// (7, 9, 'neigh_op_tnl_4')
// (7, 9, 'sp4_v_b_20')
// (7, 10, 'neigh_op_lft_4')
// (7, 10, 'sp4_v_b_9')
// (7, 10, 'sp4_v_t_44')
// (7, 11, 'neigh_op_bnl_4')
// (7, 11, 'sp4_v_b_44')
// (7, 12, 'sp4_v_b_33')
// (7, 13, 'sp4_v_b_20')
// (7, 14, 'sp4_v_b_9')

reg n305 = 0;
// (5, 9, 'neigh_op_tnr_5')
// (5, 10, 'neigh_op_rgt_5')
// (5, 11, 'neigh_op_bnr_5')
// (6, 9, 'neigh_op_top_5')
// (6, 10, 'local_g2_5')
// (6, 10, 'lutff_5/out')
// (6, 10, 'lutff_6/in_1')
// (6, 11, 'neigh_op_bot_5')
// (7, 9, 'neigh_op_tnl_5')
// (7, 10, 'neigh_op_lft_5')
// (7, 11, 'neigh_op_bnl_5')

reg n306 = 0;
// (5, 9, 'neigh_op_tnr_6')
// (5, 10, 'neigh_op_rgt_6')
// (5, 11, 'neigh_op_bnr_6')
// (6, 9, 'neigh_op_top_6')
// (6, 10, 'local_g1_6')
// (6, 10, 'lutff_0/in_1')
// (6, 10, 'lutff_6/out')
// (6, 11, 'neigh_op_bot_6')
// (7, 9, 'neigh_op_tnl_6')
// (7, 10, 'neigh_op_lft_6')
// (7, 11, 'neigh_op_bnl_6')

reg n307 = 0;
// (5, 10, 'local_g3_5')
// (5, 10, 'lutff_1/in_3')
// (5, 10, 'sp4_r_v_b_45')
// (5, 11, 'sp4_r_v_b_32')
// (5, 12, 'neigh_op_tnr_4')
// (5, 12, 'sp4_r_v_b_21')
// (5, 13, 'neigh_op_rgt_4')
// (5, 13, 'sp4_r_v_b_8')
// (5, 14, 'neigh_op_bnr_4')
// (6, 9, 'sp4_v_t_45')
// (6, 10, 'sp4_v_b_45')
// (6, 11, 'sp4_v_b_32')
// (6, 12, 'neigh_op_top_4')
// (6, 12, 'sp4_v_b_21')
// (6, 13, 'lutff_4/out')
// (6, 13, 'sp4_v_b_8')
// (6, 14, 'neigh_op_bot_4')
// (7, 12, 'neigh_op_tnl_4')
// (7, 13, 'neigh_op_lft_4')
// (7, 14, 'neigh_op_bnl_4')

reg n308 = 0;
// (5, 10, 'neigh_op_tnr_1')
// (5, 11, 'neigh_op_rgt_1')
// (5, 12, 'neigh_op_bnr_1')
// (6, 0, 'span12_vert_22')
// (6, 1, 'sp12_v_b_22')
// (6, 2, 'sp12_v_b_21')
// (6, 3, 'sp12_v_b_18')
// (6, 4, 'sp12_v_b_17')
// (6, 5, 'sp12_v_b_14')
// (6, 6, 'sp12_v_b_13')
// (6, 7, 'sp12_v_b_10')
// (6, 8, 'local_g2_1')
// (6, 8, 'lutff_7/in_0')
// (6, 8, 'sp12_v_b_9')
// (6, 9, 'sp12_v_b_6')
// (6, 10, 'neigh_op_top_1')
// (6, 10, 'sp12_v_b_5')
// (6, 11, 'local_g1_1')
// (6, 11, 'lutff_1/out')
// (6, 11, 'lutff_5/in_1')
// (6, 11, 'sp12_v_b_2')
// (6, 12, 'neigh_op_bot_1')
// (6, 12, 'sp12_v_b_1')
// (7, 10, 'neigh_op_tnl_1')
// (7, 11, 'neigh_op_lft_1')
// (7, 12, 'neigh_op_bnl_1')

reg n309 = 0;
// (5, 10, 'neigh_op_tnr_2')
// (5, 11, 'neigh_op_rgt_2')
// (5, 12, 'neigh_op_bnr_2')
// (6, 10, 'neigh_op_top_2')
// (6, 11, 'local_g1_2')
// (6, 11, 'lutff_2/out')
// (6, 11, 'lutff_4/in_1')
// (6, 11, 'lutff_7/in_2')
// (6, 12, 'neigh_op_bot_2')
// (7, 10, 'neigh_op_tnl_2')
// (7, 11, 'neigh_op_lft_2')
// (7, 12, 'neigh_op_bnl_2')

reg n310 = 0;
// (5, 10, 'neigh_op_tnr_3')
// (5, 11, 'neigh_op_rgt_3')
// (5, 12, 'neigh_op_bnr_3')
// (6, 10, 'neigh_op_top_3')
// (6, 11, 'local_g1_3')
// (6, 11, 'lutff_3/out')
// (6, 11, 'lutff_7/in_1')
// (6, 12, 'neigh_op_bot_3')
// (7, 10, 'neigh_op_tnl_3')
// (7, 11, 'neigh_op_lft_3')
// (7, 12, 'neigh_op_bnl_3')

reg n311 = 0;
// (5, 10, 'neigh_op_tnr_4')
// (5, 11, 'neigh_op_rgt_4')
// (5, 12, 'neigh_op_bnr_4')
// (6, 10, 'neigh_op_top_4')
// (6, 11, 'local_g0_4')
// (6, 11, 'lutff_0/in_2')
// (6, 11, 'lutff_1/in_1')
// (6, 11, 'lutff_4/out')
// (6, 12, 'neigh_op_bot_4')
// (7, 10, 'neigh_op_tnl_4')
// (7, 11, 'neigh_op_lft_4')
// (7, 12, 'neigh_op_bnl_4')

reg n312 = 0;
// (5, 10, 'neigh_op_tnr_5')
// (5, 11, 'neigh_op_rgt_5')
// (5, 12, 'neigh_op_bnr_5')
// (6, 10, 'neigh_op_top_5')
// (6, 11, 'local_g2_5')
// (6, 11, 'lutff_2/in_1')
// (6, 11, 'lutff_3/in_2')
// (6, 11, 'lutff_5/out')
// (6, 12, 'neigh_op_bot_5')
// (7, 10, 'neigh_op_tnl_5')
// (7, 11, 'neigh_op_lft_5')
// (7, 12, 'neigh_op_bnl_5')

reg n313 = 0;
// (5, 10, 'neigh_op_tnr_7')
// (5, 11, 'neigh_op_rgt_7')
// (5, 12, 'neigh_op_bnr_7')
// (6, 10, 'neigh_op_top_7')
// (6, 11, 'local_g0_7')
// (6, 11, 'lutff_0/in_1')
// (6, 11, 'lutff_7/out')
// (6, 12, 'neigh_op_bot_7')
// (7, 10, 'neigh_op_tnl_7')
// (7, 11, 'neigh_op_lft_7')
// (7, 12, 'neigh_op_bnl_7')

reg n314 = 0;
// (5, 11, 'neigh_op_tnr_0')
// (5, 12, 'neigh_op_rgt_0')
// (5, 13, 'neigh_op_bnr_0')
// (6, 11, 'neigh_op_top_0')
// (6, 12, 'local_g1_0')
// (6, 12, 'lutff_0/out')
// (6, 12, 'lutff_5/in_0')
// (6, 13, 'neigh_op_bot_0')
// (7, 11, 'neigh_op_tnl_0')
// (7, 12, 'neigh_op_lft_0')
// (7, 13, 'neigh_op_bnl_0')

reg n315 = 0;
// (5, 11, 'neigh_op_tnr_1')
// (5, 12, 'neigh_op_rgt_1')
// (5, 13, 'neigh_op_bnr_1')
// (6, 11, 'neigh_op_top_1')
// (6, 12, 'local_g0_1')
// (6, 12, 'lutff_1/out')
// (6, 12, 'lutff_7/in_0')
// (6, 13, 'neigh_op_bot_1')
// (7, 11, 'neigh_op_tnl_1')
// (7, 12, 'neigh_op_lft_1')
// (7, 13, 'neigh_op_bnl_1')

reg n316 = 0;
// (5, 11, 'neigh_op_tnr_2')
// (5, 12, 'neigh_op_rgt_2')
// (5, 13, 'neigh_op_bnr_2')
// (6, 11, 'neigh_op_top_2')
// (6, 12, 'lutff_2/out')
// (6, 13, 'local_g1_2')
// (6, 13, 'lutff_1/in_0')
// (6, 13, 'neigh_op_bot_2')
// (7, 11, 'neigh_op_tnl_2')
// (7, 12, 'neigh_op_lft_2')
// (7, 13, 'neigh_op_bnl_2')

reg n317 = 0;
// (5, 11, 'neigh_op_tnr_3')
// (5, 12, 'neigh_op_rgt_3')
// (5, 13, 'neigh_op_bnr_3')
// (6, 11, 'neigh_op_top_3')
// (6, 12, 'local_g1_3')
// (6, 12, 'lutff_0/in_0')
// (6, 12, 'lutff_3/out')
// (6, 13, 'neigh_op_bot_3')
// (7, 11, 'neigh_op_tnl_3')
// (7, 12, 'neigh_op_lft_3')
// (7, 13, 'neigh_op_bnl_3')

reg n318 = 0;
// (5, 11, 'neigh_op_tnr_4')
// (5, 12, 'neigh_op_rgt_4')
// (5, 13, 'neigh_op_bnr_4')
// (6, 11, 'neigh_op_top_4')
// (6, 12, 'local_g1_4')
// (6, 12, 'lutff_3/in_0')
// (6, 12, 'lutff_4/out')
// (6, 13, 'neigh_op_bot_4')
// (7, 11, 'neigh_op_tnl_4')
// (7, 12, 'neigh_op_lft_4')
// (7, 13, 'neigh_op_bnl_4')

reg n319 = 0;
// (5, 11, 'neigh_op_tnr_5')
// (5, 12, 'neigh_op_rgt_5')
// (5, 13, 'neigh_op_bnr_5')
// (6, 5, 'sp4_r_v_b_39')
// (6, 6, 'sp4_r_v_b_26')
// (6, 7, 'sp4_r_v_b_15')
// (6, 8, 'local_g1_2')
// (6, 8, 'lutff_1/in_0')
// (6, 8, 'sp4_r_v_b_2')
// (6, 9, 'sp4_r_v_b_46')
// (6, 10, 'local_g0_0')
// (6, 10, 'lutff_4/in_0')
// (6, 10, 'sp4_r_v_b_35')
// (6, 11, 'neigh_op_top_5')
// (6, 11, 'sp4_r_v_b_22')
// (6, 12, 'local_g1_5')
// (6, 12, 'lutff_4/in_0')
// (6, 12, 'lutff_5/out')
// (6, 12, 'sp4_r_v_b_11')
// (6, 13, 'neigh_op_bot_5')
// (7, 4, 'sp4_v_t_39')
// (7, 5, 'sp4_v_b_39')
// (7, 6, 'sp4_v_b_26')
// (7, 7, 'sp4_v_b_15')
// (7, 8, 'local_g1_4')
// (7, 8, 'lutff_7/in_0')
// (7, 8, 'sp4_h_r_4')
// (7, 8, 'sp4_v_b_2')
// (7, 8, 'sp4_v_t_46')
// (7, 9, 'sp4_v_b_46')
// (7, 10, 'sp4_v_b_35')
// (7, 11, 'neigh_op_tnl_5')
// (7, 11, 'sp4_v_b_22')
// (7, 12, 'neigh_op_lft_5')
// (7, 12, 'sp4_v_b_11')
// (7, 13, 'neigh_op_bnl_5')
// (8, 8, 'sp4_h_r_17')
// (9, 8, 'sp4_h_r_28')
// (10, 8, 'sp4_h_r_41')
// (11, 8, 'sp4_h_l_41')

reg n320 = 0;
// (5, 11, 'neigh_op_tnr_6')
// (5, 12, 'neigh_op_rgt_6')
// (5, 13, 'neigh_op_bnr_6')
// (6, 8, 'sp4_r_v_b_46')
// (6, 9, 'local_g0_0')
// (6, 9, 'lutff_0/in_0')
// (6, 9, 'sp4_r_v_b_35')
// (6, 10, 'sp4_r_v_b_22')
// (6, 11, 'neigh_op_top_6')
// (6, 11, 'sp4_r_v_b_11')
// (6, 12, 'local_g1_6')
// (6, 12, 'lutff_4/in_1')
// (6, 12, 'lutff_6/out')
// (6, 12, 'sp4_r_v_b_45')
// (6, 13, 'neigh_op_bot_6')
// (6, 13, 'sp4_r_v_b_32')
// (6, 14, 'sp4_r_v_b_21')
// (6, 15, 'sp4_r_v_b_8')
// (7, 7, 'sp4_v_t_46')
// (7, 8, 'sp4_v_b_46')
// (7, 9, 'sp4_v_b_35')
// (7, 10, 'sp4_v_b_22')
// (7, 11, 'neigh_op_tnl_6')
// (7, 11, 'sp4_v_b_11')
// (7, 11, 'sp4_v_t_45')
// (7, 12, 'neigh_op_lft_6')
// (7, 12, 'sp4_v_b_45')
// (7, 13, 'neigh_op_bnl_6')
// (7, 13, 'sp4_v_b_32')
// (7, 14, 'sp4_v_b_21')
// (7, 15, 'sp4_v_b_8')

reg n321 = 0;
// (5, 11, 'neigh_op_tnr_7')
// (5, 12, 'neigh_op_rgt_7')
// (5, 13, 'neigh_op_bnr_7')
// (6, 11, 'neigh_op_top_7')
// (6, 12, 'local_g1_7')
// (6, 12, 'lutff_6/in_0')
// (6, 12, 'lutff_7/out')
// (6, 13, 'neigh_op_bot_7')
// (7, 11, 'neigh_op_tnl_7')
// (7, 12, 'neigh_op_lft_7')
// (7, 13, 'neigh_op_bnl_7')

reg n322 = 0;
// (5, 12, 'neigh_op_tnr_1')
// (5, 13, 'neigh_op_rgt_1')
// (5, 14, 'neigh_op_bnr_1')
// (6, 12, 'neigh_op_top_1')
// (6, 13, 'local_g0_1')
// (6, 13, 'lutff_1/out')
// (6, 13, 'lutff_7/in_0')
// (6, 14, 'neigh_op_bot_1')
// (7, 12, 'neigh_op_tnl_1')
// (7, 13, 'neigh_op_lft_1')
// (7, 14, 'neigh_op_bnl_1')

reg n323 = 0;
// (5, 12, 'neigh_op_tnr_7')
// (5, 13, 'neigh_op_rgt_7')
// (5, 14, 'neigh_op_bnr_7')
// (6, 12, 'neigh_op_top_7')
// (6, 13, 'local_g1_7')
// (6, 13, 'lutff_4/in_0')
// (6, 13, 'lutff_7/out')
// (6, 14, 'neigh_op_bot_7')
// (7, 12, 'neigh_op_tnl_7')
// (7, 13, 'neigh_op_lft_7')
// (7, 14, 'neigh_op_bnl_7')

reg n324 = 0;
// (5, 12, 'sp12_h_r_0')
// (6, 12, 'sp12_h_r_3')
// (7, 12, 'sp12_h_r_4')
// (8, 12, 'sp12_h_r_7')
// (9, 12, 'local_g1_0')
// (9, 12, 'lutff_1/in_0')
// (9, 12, 'sp12_h_r_8')
// (10, 11, 'neigh_op_tnr_2')
// (10, 12, 'neigh_op_rgt_2')
// (10, 12, 'sp12_h_r_11')
// (10, 13, 'neigh_op_bnr_2')
// (11, 11, 'neigh_op_top_2')
// (11, 12, 'lutff_2/out')
// (11, 12, 'sp12_h_r_12')
// (11, 13, 'neigh_op_bot_2')
// (12, 11, 'neigh_op_tnl_2')
// (12, 12, 'neigh_op_lft_2')
// (12, 12, 'sp12_h_r_15')
// (12, 13, 'neigh_op_bnl_2')
// (13, 12, 'span12_horz_15')

reg n325 = 0;
// (5, 13, 'neigh_op_tnr_7')
// (5, 14, 'neigh_op_rgt_7')
// (5, 15, 'neigh_op_bnr_7')
// (6, 9, 'sp12_v_t_22')
// (6, 10, 'local_g2_6')
// (6, 10, 'lutff_5/in_1')
// (6, 10, 'sp12_v_b_22')
// (6, 11, 'sp12_v_b_21')
// (6, 12, 'sp12_v_b_18')
// (6, 13, 'neigh_op_top_7')
// (6, 13, 'sp12_v_b_17')
// (6, 14, 'lutff_7/out')
// (6, 14, 'sp12_v_b_14')
// (6, 15, 'neigh_op_bot_7')
// (6, 15, 'sp12_v_b_13')
// (6, 16, 'sp12_v_b_10')
// (6, 17, 'span12_vert_9')
// (7, 13, 'neigh_op_tnl_7')
// (7, 14, 'neigh_op_lft_7')
// (7, 15, 'neigh_op_bnl_7')

wire n326;
// (6, 0, 'logic_op_tnr_0')
// (6, 1, 'neigh_op_rgt_0')
// (6, 2, 'neigh_op_bnr_0')
// (7, 0, 'logic_op_top_0')
// (7, 1, 'local_g3_0')
// (7, 1, 'lutff_0/out')
// (7, 1, 'lutff_6/in_3')
// (7, 2, 'neigh_op_bot_0')
// (8, 0, 'logic_op_tnl_0')
// (8, 1, 'neigh_op_lft_0')
// (8, 2, 'neigh_op_bnl_0')

wire n327;
// (6, 0, 'logic_op_tnr_1')
// (6, 1, 'neigh_op_rgt_1')
// (6, 2, 'neigh_op_bnr_1')
// (7, 0, 'logic_op_top_1')
// (7, 1, 'local_g2_1')
// (7, 1, 'local_g3_1')
// (7, 1, 'lutff_1/out')
// (7, 1, 'lutff_2/in_2')
// (7, 1, 'lutff_7/in_2')
// (7, 2, 'neigh_op_bot_1')
// (8, 0, 'logic_op_tnl_1')
// (8, 1, 'neigh_op_lft_1')
// (8, 2, 'neigh_op_bnl_1')

wire n328;
// (6, 0, 'logic_op_tnr_2')
// (6, 1, 'local_g3_2')
// (6, 1, 'lutff_1/in_2')
// (6, 1, 'neigh_op_rgt_2')
// (6, 2, 'neigh_op_bnr_2')
// (7, 0, 'logic_op_top_2')
// (7, 1, 'local_g0_2')
// (7, 1, 'local_g1_2')
// (7, 1, 'lutff_2/out')
// (7, 1, 'lutff_3/in_0')
// (7, 1, 'lutff_6/in_0')
// (7, 2, 'neigh_op_bot_2')
// (8, 0, 'logic_op_tnl_2')
// (8, 1, 'neigh_op_lft_2')
// (8, 2, 'neigh_op_bnl_2')

wire n329;
// (6, 0, 'logic_op_tnr_3')
// (6, 1, 'neigh_op_rgt_3')
// (6, 2, 'neigh_op_bnr_3')
// (7, 0, 'logic_op_top_3')
// (7, 1, 'lutff_3/out')
// (7, 1, 'sp4_r_v_b_23')
// (7, 2, 'local_g1_3')
// (7, 2, 'lutff_3/in_3')
// (7, 2, 'neigh_op_bot_3')
// (7, 2, 'sp4_r_v_b_10')
// (8, 0, 'logic_op_tnl_3')
// (8, 0, 'span4_vert_23')
// (8, 1, 'neigh_op_lft_3')
// (8, 1, 'sp4_v_b_23')
// (8, 2, 'neigh_op_bnl_3')
// (8, 2, 'sp4_h_r_4')
// (8, 2, 'sp4_v_b_10')
// (9, 2, 'sp4_h_r_17')
// (10, 2, 'sp4_h_r_28')
// (11, 2, 'local_g3_1')
// (11, 2, 'lutff_7/in_3')
// (11, 2, 'sp4_h_r_41')
// (12, 2, 'sp4_h_l_41')

wire n330;
// (6, 0, 'logic_op_tnr_4')
// (6, 1, 'neigh_op_rgt_4')
// (6, 1, 'sp4_r_v_b_24')
// (6, 2, 'neigh_op_bnr_4')
// (6, 2, 'sp4_r_v_b_13')
// (6, 3, 'sp4_r_v_b_0')
// (7, 0, 'logic_op_top_4')
// (7, 0, 'span4_vert_24')
// (7, 1, 'lutff_4/out')
// (7, 1, 'sp4_v_b_24')
// (7, 2, 'neigh_op_bot_4')
// (7, 2, 'sp4_v_b_13')
// (7, 3, 'local_g0_0')
// (7, 3, 'local_g1_0')
// (7, 3, 'lutff_3/in_2')
// (7, 3, 'lutff_4/in_1')
// (7, 3, 'lutff_5/in_1')
// (7, 3, 'lutff_6/in_1')
// (7, 3, 'sp4_v_b_0')
// (8, 0, 'logic_op_tnl_4')
// (8, 1, 'neigh_op_lft_4')
// (8, 2, 'neigh_op_bnl_4')

wire n331;
// (6, 0, 'logic_op_tnr_5')
// (6, 1, 'neigh_op_rgt_5')
// (6, 2, 'neigh_op_bnr_5')
// (7, 0, 'logic_op_top_5')
// (7, 1, 'lutff_5/out')
// (7, 1, 'sp4_h_r_10')
// (7, 2, 'local_g0_5')
// (7, 2, 'lutff_6/in_1')
// (7, 2, 'neigh_op_bot_5')
// (8, 0, 'logic_op_tnl_5')
// (8, 1, 'neigh_op_lft_5')
// (8, 1, 'sp4_h_r_23')
// (8, 2, 'neigh_op_bnl_5')
// (9, 1, 'sp4_h_r_34')
// (10, 1, 'sp4_h_r_47')
// (10, 2, 'sp4_r_v_b_38')
// (10, 3, 'sp4_r_v_b_27')
// (10, 4, 'sp4_r_v_b_14')
// (10, 5, 'sp4_r_v_b_3')
// (11, 1, 'sp4_h_l_47')
// (11, 1, 'sp4_v_t_38')
// (11, 2, 'local_g2_6')
// (11, 2, 'lutff_7/in_1')
// (11, 2, 'sp4_v_b_38')
// (11, 3, 'sp4_v_b_27')
// (11, 4, 'sp4_v_b_14')
// (11, 5, 'sp4_v_b_3')

wire n332;
// (6, 0, 'logic_op_tnr_6')
// (6, 1, 'neigh_op_rgt_6')
// (6, 2, 'local_g0_6')
// (6, 2, 'lutff_5/in_3')
// (6, 2, 'neigh_op_bnr_6')
// (7, 0, 'logic_op_top_6')
// (7, 1, 'lutff_6/out')
// (7, 2, 'local_g1_6')
// (7, 2, 'lutff_6/in_3')
// (7, 2, 'neigh_op_bot_6')
// (8, 0, 'logic_op_tnl_6')
// (8, 1, 'neigh_op_lft_6')
// (8, 2, 'neigh_op_bnl_6')

wire n333;
// (6, 0, 'logic_op_tnr_7')
// (6, 1, 'local_g3_7')
// (6, 1, 'lutff_1/in_1')
// (6, 1, 'neigh_op_rgt_7')
// (6, 2, 'local_g0_7')
// (6, 2, 'local_g1_7')
// (6, 2, 'lutff_1/in_0')
// (6, 2, 'lutff_3/in_3')
// (6, 2, 'lutff_4/in_2')
// (6, 2, 'lutff_6/in_2')
// (6, 2, 'neigh_op_bnr_7')
// (7, 0, 'logic_op_top_7')
// (7, 1, 'local_g2_7')
// (7, 1, 'local_g3_7')
// (7, 1, 'lutff_4/in_0')
// (7, 1, 'lutff_5/in_0')
// (7, 1, 'lutff_7/out')
// (7, 2, 'neigh_op_bot_7')
// (8, 0, 'logic_op_tnl_7')
// (8, 1, 'neigh_op_lft_7')
// (8, 2, 'neigh_op_bnl_7')

wire n334;
// (6, 1, 'local_g3_4')
// (6, 1, 'lutff_1/in_0')
// (6, 1, 'neigh_op_tnr_4')
// (6, 2, 'local_g2_4')
// (6, 2, 'local_g3_4')
// (6, 2, 'lutff_1/in_2')
// (6, 2, 'lutff_3/in_1')
// (6, 2, 'lutff_4/in_0')
// (6, 2, 'lutff_6/in_3')
// (6, 2, 'neigh_op_rgt_4')
// (6, 3, 'neigh_op_bnr_4')
// (7, 1, 'local_g0_4')
// (7, 1, 'local_g1_4')
// (7, 1, 'lutff_3/in_1')
// (7, 1, 'lutff_4/in_2')
// (7, 1, 'lutff_5/in_1')
// (7, 1, 'lutff_6/in_1')
// (7, 1, 'neigh_op_top_4')
// (7, 2, 'lutff_4/out')
// (7, 3, 'neigh_op_bot_4')
// (8, 1, 'neigh_op_tnl_4')
// (8, 2, 'neigh_op_lft_4')
// (8, 3, 'neigh_op_bnl_4')

wire n335;
// (6, 1, 'local_g3_5')
// (6, 1, 'lutff_1/in_3')
// (6, 1, 'neigh_op_tnr_5')
// (6, 2, 'local_g2_5')
// (6, 2, 'local_g3_5')
// (6, 2, 'lutff_1/in_3')
// (6, 2, 'lutff_3/in_0')
// (6, 2, 'lutff_4/in_1')
// (6, 2, 'lutff_6/in_1')
// (6, 2, 'neigh_op_rgt_5')
// (6, 3, 'neigh_op_bnr_5')
// (7, 1, 'local_g0_5')
// (7, 1, 'local_g1_5')
// (7, 1, 'lutff_4/in_3')
// (7, 1, 'lutff_5/in_3')
// (7, 1, 'neigh_op_top_5')
// (7, 2, 'lutff_5/out')
// (7, 3, 'neigh_op_bot_5')
// (8, 1, 'neigh_op_tnl_5')
// (8, 2, 'neigh_op_lft_5')
// (8, 3, 'neigh_op_bnl_5')

wire n336;
// (6, 1, 'neigh_op_tnr_0')
// (6, 2, 'neigh_op_rgt_0')
// (6, 3, 'neigh_op_bnr_0')
// (7, 1, 'local_g0_0')
// (7, 1, 'local_g1_0')
// (7, 1, 'lutff_3/in_2')
// (7, 1, 'lutff_6/in_2')
// (7, 1, 'neigh_op_top_0')
// (7, 2, 'lutff_0/out')
// (7, 3, 'neigh_op_bot_0')
// (8, 1, 'neigh_op_tnl_0')
// (8, 2, 'neigh_op_lft_0')
// (8, 3, 'neigh_op_bnl_0')

wire n337;
// (6, 1, 'neigh_op_tnr_1')
// (6, 2, 'neigh_op_rgt_1')
// (6, 3, 'neigh_op_bnr_1')
// (7, 1, 'neigh_op_top_1')
// (7, 2, 'local_g0_1')
// (7, 2, 'local_g1_1')
// (7, 2, 'lutff_0/in_1')
// (7, 2, 'lutff_1/out')
// (7, 2, 'lutff_4/in_2')
// (7, 2, 'lutff_5/in_2')
// (7, 3, 'neigh_op_bot_1')
// (8, 1, 'neigh_op_tnl_1')
// (8, 2, 'neigh_op_lft_1')
// (8, 3, 'neigh_op_bnl_1')

wire n338;
// (6, 1, 'neigh_op_tnr_2')
// (6, 1, 'sp4_r_v_b_17')
// (6, 2, 'neigh_op_rgt_2')
// (6, 2, 'sp4_r_v_b_4')
// (6, 3, 'neigh_op_bnr_2')
// (7, 0, 'span4_vert_17')
// (7, 1, 'local_g0_1')
// (7, 1, 'local_g1_1')
// (7, 1, 'lutff_2/in_1')
// (7, 1, 'lutff_7/in_1')
// (7, 1, 'neigh_op_top_2')
// (7, 1, 'sp4_v_b_17')
// (7, 2, 'lutff_2/out')
// (7, 2, 'sp4_v_b_4')
// (7, 3, 'neigh_op_bot_2')
// (8, 1, 'neigh_op_tnl_2')
// (8, 2, 'neigh_op_lft_2')
// (8, 3, 'neigh_op_bnl_2')

wire n339;
// (6, 1, 'neigh_op_tnr_3')
// (6, 2, 'neigh_op_rgt_3')
// (6, 3, 'neigh_op_bnr_3')
// (7, 1, 'neigh_op_top_3')
// (7, 2, 'lutff_3/out')
// (7, 3, 'local_g0_3')
// (7, 3, 'lutff_1/in_2')
// (7, 3, 'neigh_op_bot_3')
// (8, 1, 'neigh_op_tnl_3')
// (8, 2, 'neigh_op_lft_3')
// (8, 3, 'neigh_op_bnl_3')

wire n340;
// (6, 1, 'neigh_op_tnr_7')
// (6, 2, 'neigh_op_rgt_7')
// (6, 3, 'neigh_op_bnr_7')
// (7, 1, 'local_g0_7')
// (7, 1, 'local_g1_7')
// (7, 1, 'lutff_2/in_3')
// (7, 1, 'lutff_7/in_3')
// (7, 1, 'neigh_op_top_7')
// (7, 2, 'lutff_7/out')
// (7, 3, 'neigh_op_bot_7')
// (8, 1, 'neigh_op_tnl_7')
// (8, 2, 'local_g1_7')
// (8, 2, 'lutff_2/in_2')
// (8, 2, 'lutff_4/in_2')
// (8, 2, 'neigh_op_lft_7')
// (8, 3, 'neigh_op_bnl_7')

wire n341;
// (6, 1, 'sp4_r_v_b_19')
// (6, 2, 'sp4_r_v_b_6')
// (7, 0, 'span4_vert_19')
// (7, 1, 'local_g2_6')
// (7, 1, 'lutff_0/in_2')
// (7, 1, 'lutff_1/in_1')
// (7, 1, 'neigh_op_tnr_6')
// (7, 1, 'sp4_v_b_19')
// (7, 2, 'local_g0_6')
// (7, 2, 'lutff_6/in_0')
// (7, 2, 'neigh_op_rgt_6')
// (7, 2, 'sp4_h_r_1')
// (7, 2, 'sp4_v_b_6')
// (7, 3, 'neigh_op_bnr_6')
// (8, 1, 'neigh_op_top_6')
// (8, 2, 'local_g3_6')
// (8, 2, 'lutff_0/in_1')
// (8, 2, 'lutff_6/out')
// (8, 2, 'sp4_h_r_12')
// (8, 3, 'neigh_op_bot_6')
// (9, 1, 'neigh_op_tnl_6')
// (9, 2, 'neigh_op_lft_6')
// (9, 2, 'sp4_h_r_25')
// (9, 3, 'neigh_op_bnl_6')
// (10, 2, 'sp4_h_r_36')
// (11, 2, 'sp4_h_l_36')

wire n342;
// (6, 1, 'sp4_r_v_b_27')
// (6, 1, 'sp4_r_v_b_32')
// (6, 2, 'local_g2_6')
// (6, 2, 'lutff_7/in_3')
// (6, 2, 'sp4_r_v_b_14')
// (6, 2, 'sp4_r_v_b_21')
// (6, 3, 'local_g2_0')
// (6, 3, 'lutff_3/in_1')
// (6, 3, 'sp4_r_v_b_3')
// (6, 3, 'sp4_r_v_b_8')
// (7, 0, 'span4_vert_27')
// (7, 0, 'span4_vert_32')
// (7, 1, 'sp4_r_v_b_38')
// (7, 1, 'sp4_v_b_27')
// (7, 1, 'sp4_v_b_32')
// (7, 2, 'neigh_op_tnr_7')
// (7, 2, 'sp4_r_v_b_27')
// (7, 2, 'sp4_v_b_14')
// (7, 2, 'sp4_v_b_21')
// (7, 3, 'neigh_op_rgt_7')
// (7, 3, 'sp4_h_r_3')
// (7, 3, 'sp4_r_v_b_14')
// (7, 3, 'sp4_v_b_3')
// (7, 3, 'sp4_v_b_8')
// (7, 4, 'neigh_op_bnr_7')
// (7, 4, 'sp4_r_v_b_3')
// (8, 0, 'span4_vert_38')
// (8, 1, 'sp4_v_b_38')
// (8, 2, 'local_g2_3')
// (8, 2, 'lutff_1/in_0')
// (8, 2, 'lutff_7/in_0')
// (8, 2, 'neigh_op_top_7')
// (8, 2, 'sp4_v_b_27')
// (8, 3, 'lutff_7/out')
// (8, 3, 'sp4_h_r_14')
// (8, 3, 'sp4_v_b_14')
// (8, 4, 'neigh_op_bot_7')
// (8, 4, 'sp4_v_b_3')
// (9, 2, 'neigh_op_tnl_7')
// (9, 3, 'neigh_op_lft_7')
// (9, 3, 'sp4_h_r_27')
// (9, 4, 'neigh_op_bnl_7')
// (10, 3, 'sp4_h_r_38')
// (11, 3, 'sp4_h_l_38')

reg n343 = 0;
// (6, 1, 'sp4_r_v_b_29')
// (6, 2, 'sp4_r_v_b_16')
// (6, 3, 'sp4_r_v_b_5')
// (6, 4, 'sp4_r_v_b_39')
// (6, 5, 'sp4_r_v_b_26')
// (6, 6, 'sp4_r_v_b_15')
// (6, 7, 'sp4_r_v_b_2')
// (6, 8, 'sp4_r_v_b_43')
// (6, 9, 'sp4_r_v_b_30')
// (6, 10, 'sp4_r_v_b_19')
// (6, 11, 'sp4_r_v_b_6')
// (7, 0, 'span4_vert_29')
// (7, 1, 'sp4_v_b_29')
// (7, 2, 'sp4_v_b_16')
// (7, 3, 'local_g0_5')
// (7, 3, 'lutff_0/in_3')
// (7, 3, 'sp4_v_b_5')
// (7, 3, 'sp4_v_t_39')
// (7, 4, 'sp4_v_b_39')
// (7, 5, 'sp4_v_b_26')
// (7, 6, 'sp4_v_b_15')
// (7, 7, 'sp4_v_b_2')
// (7, 7, 'sp4_v_t_43')
// (7, 8, 'sp4_v_b_43')
// (7, 9, 'sp4_v_b_30')
// (7, 10, 'sp4_v_b_19')
// (7, 11, 'sp4_h_r_6')
// (7, 11, 'sp4_v_b_6')
// (8, 10, 'neigh_op_tnr_7')
// (8, 11, 'neigh_op_rgt_7')
// (8, 11, 'sp4_h_r_19')
// (8, 12, 'neigh_op_bnr_7')
// (9, 10, 'neigh_op_top_7')
// (9, 11, 'local_g1_7')
// (9, 11, 'lutff_1/in_1')
// (9, 11, 'lutff_7/out')
// (9, 11, 'sp4_h_r_30')
// (9, 12, 'neigh_op_bot_7')
// (10, 10, 'neigh_op_tnl_7')
// (10, 11, 'neigh_op_lft_7')
// (10, 11, 'sp4_h_r_43')
// (10, 12, 'neigh_op_bnl_7')
// (11, 11, 'sp4_h_l_43')

wire n344;
// (6, 1, 'sp4_r_v_b_34')
// (6, 2, 'local_g3_7')
// (6, 2, 'lutff_2/in_2')
// (6, 2, 'neigh_op_tnr_5')
// (6, 2, 'sp4_r_v_b_23')
// (6, 3, 'neigh_op_rgt_5')
// (6, 3, 'sp4_r_v_b_10')
// (6, 4, 'neigh_op_bnr_5')
// (7, 0, 'span4_vert_34')
// (7, 1, 'sp4_v_b_34')
// (7, 2, 'local_g0_7')
// (7, 2, 'lutff_3/in_2')
// (7, 2, 'neigh_op_top_5')
// (7, 2, 'sp4_v_b_23')
// (7, 3, 'lutff_5/out')
// (7, 3, 'sp4_v_b_10')
// (7, 4, 'neigh_op_bot_5')
// (8, 2, 'neigh_op_tnl_5')
// (8, 3, 'neigh_op_lft_5')
// (8, 4, 'neigh_op_bnl_5')

wire n345;
// (6, 2, 'neigh_op_tnr_0')
// (6, 3, 'neigh_op_rgt_0')
// (6, 4, 'neigh_op_bnr_0')
// (6, 11, 'sp4_h_r_1')
// (7, 0, 'span12_vert_20')
// (7, 1, 'sp12_v_b_20')
// (7, 2, 'neigh_op_top_0')
// (7, 2, 'sp12_v_b_19')
// (7, 3, 'lutff_0/out')
// (7, 3, 'sp12_v_b_16')
// (7, 4, 'neigh_op_bot_0')
// (7, 4, 'sp12_v_b_15')
// (7, 5, 'sp12_v_b_12')
// (7, 6, 'sp12_v_b_11')
// (7, 7, 'sp12_v_b_8')
// (7, 8, 'sp12_v_b_7')
// (7, 9, 'sp12_v_b_4')
// (7, 10, 'sp12_v_b_3')
// (7, 11, 'local_g1_4')
// (7, 11, 'lutff_7/in_2')
// (7, 11, 'sp12_h_r_0')
// (7, 11, 'sp12_v_b_0')
// (7, 11, 'sp4_h_r_12')
// (8, 2, 'neigh_op_tnl_0')
// (8, 3, 'neigh_op_lft_0')
// (8, 4, 'neigh_op_bnl_0')
// (8, 11, 'sp12_h_r_3')
// (8, 11, 'sp4_h_r_25')
// (8, 11, 'sp4_h_r_3')
// (9, 11, 'sp12_h_r_4')
// (9, 11, 'sp4_h_r_14')
// (9, 11, 'sp4_h_r_36')
// (10, 11, 'sp12_h_r_7')
// (10, 11, 'sp4_h_l_36')
// (10, 11, 'sp4_h_r_27')
// (11, 8, 'local_g2_6')
// (11, 8, 'lutff_2/in_0')
// (11, 8, 'sp4_r_v_b_38')
// (11, 9, 'sp4_r_v_b_27')
// (11, 10, 'sp4_r_v_b_14')
// (11, 11, 'local_g1_0')
// (11, 11, 'lutff_5/in_2')
// (11, 11, 'sp12_h_r_8')
// (11, 11, 'sp4_h_r_38')
// (11, 11, 'sp4_r_v_b_3')
// (12, 7, 'sp4_v_t_38')
// (12, 8, 'sp4_v_b_38')
// (12, 9, 'sp4_v_b_27')
// (12, 10, 'sp4_v_b_14')
// (12, 11, 'sp12_h_r_11')
// (12, 11, 'sp4_h_l_38')
// (12, 11, 'sp4_v_b_3')
// (13, 11, 'span12_horz_11')

wire n346;
// (6, 2, 'neigh_op_tnr_1')
// (6, 3, 'neigh_op_rgt_1')
// (6, 4, 'neigh_op_bnr_1')
// (7, 2, 'neigh_op_top_1')
// (7, 3, 'lutff_1/out')
// (7, 4, 'local_g0_1')
// (7, 4, 'lutff_0/in_1')
// (7, 4, 'neigh_op_bot_1')
// (8, 2, 'neigh_op_tnl_1')
// (8, 3, 'neigh_op_lft_1')
// (8, 4, 'neigh_op_bnl_1')

wire n347;
// (6, 2, 'neigh_op_tnr_3')
// (6, 3, 'local_g2_3')
// (6, 3, 'local_g3_3')
// (6, 3, 'lutff_1/in_2')
// (6, 3, 'lutff_2/in_2')
// (6, 3, 'lutff_7/in_0')
// (6, 3, 'neigh_op_rgt_3')
// (6, 4, 'neigh_op_bnr_3')
// (7, 2, 'neigh_op_top_3')
// (7, 3, 'lutff_3/out')
// (7, 4, 'neigh_op_bot_3')
// (8, 2, 'neigh_op_tnl_3')
// (8, 3, 'neigh_op_lft_3')
// (8, 4, 'neigh_op_bnl_3')

wire n348;
// (6, 2, 'neigh_op_tnr_4')
// (6, 3, 'local_g2_4')
// (6, 3, 'local_g3_4')
// (6, 3, 'lutff_5/in_2')
// (6, 3, 'lutff_7/in_1')
// (6, 3, 'neigh_op_rgt_4')
// (6, 4, 'neigh_op_bnr_4')
// (7, 2, 'local_g0_4')
// (7, 2, 'lutff_6/in_2')
// (7, 2, 'neigh_op_top_4')
// (7, 3, 'lutff_4/out')
// (7, 4, 'neigh_op_bot_4')
// (8, 2, 'neigh_op_tnl_4')
// (8, 3, 'neigh_op_lft_4')
// (8, 4, 'neigh_op_bnl_4')

wire n349;
// (6, 2, 'neigh_op_tnr_7')
// (6, 3, 'neigh_op_rgt_7')
// (6, 4, 'neigh_op_bnr_7')
// (6, 8, 'sp4_r_v_b_36')
// (6, 9, 'sp4_r_v_b_25')
// (6, 10, 'sp4_r_v_b_12')
// (6, 11, 'sp4_r_v_b_1')
// (7, 0, 'span12_vert_18')
// (7, 1, 'sp12_v_b_18')
// (7, 2, 'neigh_op_top_7')
// (7, 2, 'sp12_v_b_17')
// (7, 3, 'lutff_7/out')
// (7, 3, 'sp12_v_b_14')
// (7, 4, 'neigh_op_bot_7')
// (7, 4, 'sp12_v_b_13')
// (7, 5, 'sp12_v_b_10')
// (7, 6, 'sp12_v_b_9')
// (7, 7, 'sp12_v_b_6')
// (7, 7, 'sp4_v_t_36')
// (7, 8, 'sp12_v_b_5')
// (7, 8, 'sp4_v_b_36')
// (7, 9, 'sp12_v_b_2')
// (7, 9, 'sp4_v_b_25')
// (7, 10, 'sp12_v_b_1')
// (7, 10, 'sp4_v_b_12')
// (7, 11, 'local_g0_1')
// (7, 11, 'lutff_5/in_2')
// (7, 11, 'sp4_v_b_1')
// (8, 2, 'neigh_op_tnl_7')
// (8, 3, 'neigh_op_lft_7')
// (8, 4, 'neigh_op_bnl_7')

reg n350 = 0;
// (6, 3, 'neigh_op_tnr_1')
// (6, 4, 'neigh_op_rgt_1')
// (6, 5, 'neigh_op_bnr_1')
// (7, 2, 'sp4_r_v_b_43')
// (7, 3, 'neigh_op_top_1')
// (7, 3, 'sp4_r_v_b_30')
// (7, 4, 'lutff_1/out')
// (7, 4, 'sp4_r_v_b_19')
// (7, 5, 'neigh_op_bot_1')
// (7, 5, 'sp4_r_v_b_6')
// (8, 1, 'sp4_v_t_43')
// (8, 2, 'sp4_v_b_43')
// (8, 3, 'neigh_op_tnl_1')
// (8, 3, 'sp4_v_b_30')
// (8, 4, 'neigh_op_lft_1')
// (8, 4, 'sp4_v_b_19')
// (8, 5, 'neigh_op_bnl_1')
// (8, 5, 'sp4_h_r_6')
// (8, 5, 'sp4_v_b_6')
// (9, 5, 'local_g0_3')
// (9, 5, 'lutff_7/in_0')
// (9, 5, 'sp4_h_r_19')
// (10, 5, 'sp4_h_r_30')
// (11, 5, 'sp4_h_r_43')
// (12, 5, 'sp4_h_l_43')

wire n351;
// (6, 4, 'local_g2_0')
// (6, 4, 'local_g3_0')
// (6, 4, 'lutff_0/in_0')
// (6, 4, 'lutff_2/in_0')
// (6, 4, 'lutff_3/in_2')
// (6, 4, 'lutff_7/in_0')
// (6, 4, 'neigh_op_tnr_0')
// (6, 5, 'local_g2_0')
// (6, 5, 'local_g3_0')
// (6, 5, 'lutff_4/in_1')
// (6, 5, 'lutff_5/in_2')
// (6, 5, 'lutff_6/in_2')
// (6, 5, 'lutff_7/in_1')
// (6, 5, 'neigh_op_rgt_0')
// (6, 6, 'neigh_op_bnr_0')
// (7, 4, 'neigh_op_top_0')
// (7, 5, 'lutff_0/out')
// (7, 6, 'neigh_op_bot_0')
// (8, 4, 'neigh_op_tnl_0')
// (8, 5, 'neigh_op_lft_0')
// (8, 6, 'neigh_op_bnl_0')

wire n352;
// (6, 4, 'local_g2_2')
// (6, 4, 'local_g3_2')
// (6, 4, 'lutff_0/in_3')
// (6, 4, 'lutff_2/in_1')
// (6, 4, 'lutff_3/in_0')
// (6, 4, 'lutff_7/in_1')
// (6, 4, 'neigh_op_tnr_2')
// (6, 5, 'local_g2_2')
// (6, 5, 'local_g3_2')
// (6, 5, 'lutff_4/in_3')
// (6, 5, 'lutff_5/in_1')
// (6, 5, 'lutff_6/in_3')
// (6, 5, 'lutff_7/in_3')
// (6, 5, 'neigh_op_rgt_2')
// (6, 6, 'neigh_op_bnr_2')
// (7, 4, 'neigh_op_top_2')
// (7, 5, 'lutff_2/out')
// (7, 6, 'neigh_op_bot_2')
// (8, 4, 'neigh_op_tnl_2')
// (8, 5, 'neigh_op_lft_2')
// (8, 6, 'neigh_op_bnl_2')

wire n353;
// (6, 4, 'local_g2_3')
// (6, 4, 'local_g3_3')
// (6, 4, 'lutff_0/in_2')
// (6, 4, 'lutff_2/in_3')
// (6, 4, 'lutff_3/in_3')
// (6, 4, 'lutff_7/in_2')
// (6, 4, 'neigh_op_tnr_3')
// (6, 5, 'local_g2_3')
// (6, 5, 'local_g3_3')
// (6, 5, 'lutff_4/in_0')
// (6, 5, 'lutff_5/in_0')
// (6, 5, 'lutff_6/in_0')
// (6, 5, 'lutff_7/in_0')
// (6, 5, 'neigh_op_rgt_3')
// (6, 6, 'neigh_op_bnr_3')
// (7, 4, 'neigh_op_top_3')
// (7, 5, 'lutff_3/out')
// (7, 6, 'neigh_op_bot_3')
// (8, 4, 'neigh_op_tnl_3')
// (8, 5, 'neigh_op_lft_3')
// (8, 6, 'neigh_op_bnl_3')

wire n354;
// (6, 4, 'local_g2_7')
// (6, 4, 'local_g3_7')
// (6, 4, 'lutff_0/in_1')
// (6, 4, 'lutff_2/in_2')
// (6, 4, 'lutff_3/in_1')
// (6, 4, 'lutff_7/in_3')
// (6, 4, 'neigh_op_tnr_7')
// (6, 5, 'local_g2_7')
// (6, 5, 'local_g3_7')
// (6, 5, 'lutff_4/in_2')
// (6, 5, 'lutff_5/in_3')
// (6, 5, 'lutff_6/in_1')
// (6, 5, 'lutff_7/in_2')
// (6, 5, 'neigh_op_rgt_7')
// (6, 6, 'neigh_op_bnr_7')
// (7, 4, 'neigh_op_top_7')
// (7, 5, 'lutff_7/out')
// (7, 6, 'neigh_op_bot_7')
// (8, 4, 'neigh_op_tnl_7')
// (8, 5, 'neigh_op_lft_7')
// (8, 6, 'neigh_op_bnl_7')

wire n355;
// (6, 4, 'neigh_op_tnr_4')
// (6, 5, 'neigh_op_rgt_4')
// (6, 6, 'neigh_op_bnr_4')
// (7, 4, 'neigh_op_top_4')
// (7, 4, 'sp4_r_v_b_36')
// (7, 5, 'local_g1_1')
// (7, 5, 'local_g1_4')
// (7, 5, 'lutff_2/in_1')
// (7, 5, 'lutff_3/in_3')
// (7, 5, 'lutff_4/out')
// (7, 5, 'sp4_r_v_b_25')
// (7, 6, 'neigh_op_bot_4')
// (7, 6, 'sp4_r_v_b_12')
// (7, 7, 'sp4_r_v_b_1')
// (8, 3, 'sp4_v_t_36')
// (8, 4, 'neigh_op_tnl_4')
// (8, 4, 'sp4_v_b_36')
// (8, 5, 'neigh_op_lft_4')
// (8, 5, 'sp4_v_b_25')
// (8, 6, 'neigh_op_bnl_4')
// (8, 6, 'sp4_v_b_12')
// (8, 7, 'sp4_v_b_1')

wire n356;
// (6, 4, 'neigh_op_tnr_5')
// (6, 5, 'neigh_op_rgt_5')
// (6, 6, 'neigh_op_bnr_5')
// (7, 4, 'neigh_op_top_5')
// (7, 5, 'local_g0_5')
// (7, 5, 'local_g3_5')
// (7, 5, 'lutff_2/in_2')
// (7, 5, 'lutff_5/out')
// (7, 5, 'lutff_7/in_2')
// (7, 6, 'neigh_op_bot_5')
// (8, 4, 'neigh_op_tnl_5')
// (8, 5, 'neigh_op_lft_5')
// (8, 6, 'neigh_op_bnl_5')

wire n357;
// (6, 4, 'neigh_op_tnr_6')
// (6, 5, 'neigh_op_rgt_6')
// (6, 6, 'neigh_op_bnr_6')
// (7, 4, 'neigh_op_top_6')
// (7, 5, 'local_g2_6')
// (7, 5, 'lutff_0/in_2')
// (7, 5, 'lutff_6/out')
// (7, 5, 'lutff_7/in_1')
// (7, 6, 'neigh_op_bot_6')
// (8, 4, 'neigh_op_tnl_6')
// (8, 5, 'neigh_op_lft_6')
// (8, 6, 'neigh_op_bnl_6')

wire n358;
// (6, 4, 'sp4_h_r_10')
// (7, 1, 'sp4_r_v_b_42')
// (7, 2, 'sp4_r_v_b_31')
// (7, 3, 'neigh_op_tnr_1')
// (7, 3, 'sp4_r_v_b_18')
// (7, 4, 'neigh_op_rgt_1')
// (7, 4, 'sp4_h_r_23')
// (7, 4, 'sp4_r_v_b_7')
// (7, 5, 'neigh_op_bnr_1')
// (8, 0, 'span4_vert_42')
// (8, 1, 'sp4_v_b_42')
// (8, 2, 'sp4_v_b_31')
// (8, 3, 'neigh_op_top_1')
// (8, 3, 'sp4_v_b_18')
// (8, 4, 'local_g0_7')
// (8, 4, 'local_g2_2')
// (8, 4, 'lutff_1/out')
// (8, 4, 'lutff_6/in_3')
// (8, 4, 'lutff_7/in_3')
// (8, 4, 'sp4_h_r_2')
// (8, 4, 'sp4_h_r_34')
// (8, 4, 'sp4_v_b_7')
// (8, 5, 'neigh_op_bot_1')
// (9, 3, 'neigh_op_tnl_1')
// (9, 4, 'neigh_op_lft_1')
// (9, 4, 'sp4_h_r_15')
// (9, 4, 'sp4_h_r_47')
// (9, 5, 'neigh_op_bnl_1')
// (10, 4, 'sp4_h_l_47')
// (10, 4, 'sp4_h_r_26')
// (11, 4, 'sp4_h_r_39')
// (12, 4, 'sp4_h_l_39')

wire n359;
// (6, 4, 'sp4_r_v_b_37')
// (6, 5, 'sp4_r_v_b_24')
// (6, 6, 'neigh_op_tnr_0')
// (6, 6, 'sp4_r_v_b_13')
// (6, 7, 'neigh_op_rgt_0')
// (6, 7, 'sp4_r_v_b_0')
// (6, 8, 'neigh_op_bnr_0')
// (7, 3, 'sp4_v_t_37')
// (7, 4, 'sp4_v_b_37')
// (7, 5, 'sp4_v_b_24')
// (7, 6, 'local_g0_0')
// (7, 6, 'local_g0_5')
// (7, 6, 'lutff_4/in_2')
// (7, 6, 'lutff_5/in_2')
// (7, 6, 'neigh_op_top_0')
// (7, 6, 'sp4_v_b_13')
// (7, 7, 'lutff_0/out')
// (7, 7, 'sp4_v_b_0')
// (7, 8, 'neigh_op_bot_0')
// (8, 6, 'neigh_op_tnl_0')
// (8, 7, 'neigh_op_lft_0')
// (8, 8, 'neigh_op_bnl_0')

wire n360;
// (6, 4, 'sp4_r_v_b_43')
// (6, 5, 'sp4_r_v_b_30')
// (6, 6, 'sp4_r_v_b_19')
// (6, 7, 'sp4_r_v_b_6')
// (6, 10, 'neigh_op_tnr_2')
// (6, 11, 'neigh_op_rgt_2')
// (6, 12, 'neigh_op_bnr_2')
// (7, 1, 'sp12_v_t_23')
// (7, 2, 'sp12_v_b_23')
// (7, 3, 'sp12_v_b_20')
// (7, 3, 'sp4_v_t_43')
// (7, 4, 'sp12_v_b_19')
// (7, 4, 'sp4_v_b_43')
// (7, 5, 'sp12_v_b_16')
// (7, 5, 'sp4_v_b_30')
// (7, 6, 'local_g1_3')
// (7, 6, 'local_g2_7')
// (7, 6, 'lutff_2/in_3')
// (7, 6, 'lutff_3/in_1')
// (7, 6, 'sp12_v_b_15')
// (7, 6, 'sp4_v_b_19')
// (7, 7, 'local_g2_4')
// (7, 7, 'lutff_0/in_2')
// (7, 7, 'sp12_v_b_12')
// (7, 7, 'sp4_v_b_6')
// (7, 8, 'sp12_v_b_11')
// (7, 9, 'sp12_v_b_8')
// (7, 10, 'neigh_op_top_2')
// (7, 10, 'sp12_v_b_7')
// (7, 11, 'lutff_2/out')
// (7, 11, 'sp12_v_b_4')
// (7, 12, 'neigh_op_bot_2')
// (7, 12, 'sp12_v_b_3')
// (7, 13, 'sp12_v_b_0')
// (8, 10, 'neigh_op_tnl_2')
// (8, 11, 'neigh_op_lft_2')
// (8, 12, 'neigh_op_bnl_2')

wire n361;
// (6, 5, 'local_g2_4')
// (6, 5, 'local_g3_4')
// (6, 5, 'lutff_0/in_3')
// (6, 5, 'lutff_3/in_3')
// (6, 5, 'neigh_op_tnr_4')
// (6, 6, 'neigh_op_rgt_4')
// (6, 7, 'neigh_op_bnr_4')
// (7, 5, 'local_g0_4')
// (7, 5, 'lutff_0/in_0')
// (7, 5, 'lutff_3/in_1')
// (7, 5, 'lutff_5/in_3')
// (7, 5, 'neigh_op_top_4')
// (7, 6, 'lutff_4/out')
// (7, 7, 'neigh_op_bot_4')
// (8, 5, 'neigh_op_tnl_4')
// (8, 6, 'neigh_op_lft_4')
// (8, 7, 'neigh_op_bnl_4')

wire n362;
// (6, 5, 'neigh_op_tnr_1')
// (6, 6, 'neigh_op_rgt_1')
// (6, 7, 'neigh_op_bnr_1')
// (7, 4, 'sp4_r_v_b_43')
// (7, 5, 'local_g0_6')
// (7, 5, 'lutff_7/in_3')
// (7, 5, 'neigh_op_top_1')
// (7, 5, 'sp4_r_v_b_30')
// (7, 6, 'lutff_1/out')
// (7, 6, 'sp4_r_v_b_19')
// (7, 7, 'neigh_op_bot_1')
// (7, 7, 'sp4_r_v_b_6')
// (8, 3, 'sp4_v_t_43')
// (8, 4, 'sp4_v_b_43')
// (8, 5, 'neigh_op_tnl_1')
// (8, 5, 'sp4_v_b_30')
// (8, 6, 'neigh_op_lft_1')
// (8, 6, 'sp4_v_b_19')
// (8, 7, 'neigh_op_bnl_1')
// (8, 7, 'sp4_v_b_6')

wire n363;
// (6, 5, 'neigh_op_tnr_3')
// (6, 6, 'neigh_op_rgt_3')
// (6, 7, 'neigh_op_bnr_3')
// (7, 5, 'local_g0_3')
// (7, 5, 'lutff_0/in_3')
// (7, 5, 'neigh_op_top_3')
// (7, 6, 'lutff_3/out')
// (7, 7, 'neigh_op_bot_3')
// (8, 5, 'neigh_op_tnl_3')
// (8, 6, 'neigh_op_lft_3')
// (8, 7, 'neigh_op_bnl_3')

wire n364;
// (6, 5, 'neigh_op_tnr_6')
// (6, 6, 'neigh_op_rgt_6')
// (6, 7, 'neigh_op_bnr_6')
// (7, 5, 'local_g1_6')
// (7, 5, 'lutff_3/in_2')
// (7, 5, 'neigh_op_top_6')
// (7, 6, 'lutff_6/out')
// (7, 7, 'neigh_op_bot_6')
// (8, 5, 'neigh_op_tnl_6')
// (8, 6, 'neigh_op_lft_6')
// (8, 7, 'neigh_op_bnl_6')

reg n365 = 0;
// (6, 5, 'neigh_op_tnr_7')
// (6, 6, 'neigh_op_rgt_7')
// (6, 6, 'sp4_h_r_3')
// (6, 7, 'neigh_op_bnr_7')
// (7, 5, 'neigh_op_top_7')
// (7, 6, 'lutff_7/out')
// (7, 6, 'sp4_h_r_14')
// (7, 7, 'neigh_op_bot_7')
// (8, 5, 'neigh_op_tnl_7')
// (8, 6, 'neigh_op_lft_7')
// (8, 6, 'sp4_h_r_27')
// (8, 7, 'neigh_op_bnl_7')
// (9, 6, 'local_g2_6')
// (9, 6, 'lutff_4/in_0')
// (9, 6, 'sp4_h_r_38')
// (10, 6, 'sp4_h_l_38')

reg n366 = 0;
// (6, 6, 'neigh_op_tnr_1')
// (6, 7, 'neigh_op_rgt_1')
// (6, 8, 'neigh_op_bnr_1')
// (7, 6, 'neigh_op_top_1')
// (7, 7, 'local_g0_1')
// (7, 7, 'lutff_1/out')
// (7, 7, 'lutff_5/in_0')
// (7, 8, 'neigh_op_bot_1')
// (8, 6, 'neigh_op_tnl_1')
// (8, 7, 'neigh_op_lft_1')
// (8, 8, 'neigh_op_bnl_1')

reg n367 = 0;
// (6, 6, 'neigh_op_tnr_2')
// (6, 7, 'neigh_op_rgt_2')
// (6, 8, 'neigh_op_bnr_2')
// (7, 6, 'neigh_op_top_2')
// (7, 7, 'local_g0_2')
// (7, 7, 'lutff_2/out')
// (7, 7, 'lutff_4/in_0')
// (7, 8, 'neigh_op_bot_2')
// (8, 6, 'neigh_op_tnl_2')
// (8, 7, 'local_g0_2')
// (8, 7, 'lutff_3/in_3')
// (8, 7, 'neigh_op_lft_2')
// (8, 8, 'neigh_op_bnl_2')

reg n368 = 0;
// (6, 6, 'neigh_op_tnr_3')
// (6, 7, 'neigh_op_rgt_3')
// (6, 8, 'neigh_op_bnr_3')
// (7, 6, 'neigh_op_top_3')
// (7, 7, 'local_g0_3')
// (7, 7, 'lutff_1/in_0')
// (7, 7, 'lutff_3/out')
// (7, 8, 'neigh_op_bot_3')
// (8, 6, 'neigh_op_tnl_3')
// (8, 7, 'neigh_op_lft_3')
// (8, 8, 'neigh_op_bnl_3')

reg n369 = 0;
// (6, 6, 'neigh_op_tnr_4')
// (6, 6, 'sp4_r_v_b_37')
// (6, 7, 'neigh_op_rgt_4')
// (6, 7, 'sp4_r_v_b_24')
// (6, 8, 'neigh_op_bnr_4')
// (6, 8, 'sp4_r_v_b_13')
// (6, 9, 'sp4_r_v_b_0')
// (6, 10, 'sp4_r_v_b_38')
// (6, 11, 'sp4_r_v_b_27')
// (6, 12, 'sp4_r_v_b_14')
// (6, 13, 'sp4_r_v_b_3')
// (7, 4, 'sp4_r_v_b_44')
// (7, 5, 'sp4_r_v_b_33')
// (7, 5, 'sp4_v_t_37')
// (7, 6, 'neigh_op_top_4')
// (7, 6, 'sp4_r_v_b_20')
// (7, 6, 'sp4_v_b_37')
// (7, 7, 'lutff_4/out')
// (7, 7, 'sp4_r_v_b_9')
// (7, 7, 'sp4_v_b_24')
// (7, 8, 'neigh_op_bot_4')
// (7, 8, 'sp4_r_v_b_37')
// (7, 8, 'sp4_v_b_13')
// (7, 9, 'local_g1_0')
// (7, 9, 'lutff_1/in_0')
// (7, 9, 'sp4_r_v_b_24')
// (7, 9, 'sp4_v_b_0')
// (7, 9, 'sp4_v_t_38')
// (7, 10, 'sp4_r_v_b_13')
// (7, 10, 'sp4_v_b_38')
// (7, 11, 'local_g3_3')
// (7, 11, 'lutff_2/in_2')
// (7, 11, 'sp4_r_v_b_0')
// (7, 11, 'sp4_v_b_27')
// (7, 12, 'sp4_v_b_14')
// (7, 13, 'sp4_v_b_3')
// (8, 3, 'sp4_v_t_44')
// (8, 4, 'sp4_v_b_44')
// (8, 5, 'sp4_v_b_33')
// (8, 6, 'neigh_op_tnl_4')
// (8, 6, 'sp4_v_b_20')
// (8, 7, 'local_g1_4')
// (8, 7, 'lutff_7/in_0')
// (8, 7, 'neigh_op_lft_4')
// (8, 7, 'sp4_v_b_9')
// (8, 7, 'sp4_v_t_37')
// (8, 8, 'neigh_op_bnl_4')
// (8, 8, 'sp4_v_b_37')
// (8, 9, 'sp4_v_b_24')
// (8, 10, 'sp4_v_b_13')
// (8, 11, 'local_g1_0')
// (8, 11, 'lutff_3/in_2')
// (8, 11, 'sp4_v_b_0')

reg n370 = 0;
// (6, 6, 'neigh_op_tnr_6')
// (6, 7, 'neigh_op_rgt_6')
// (6, 8, 'neigh_op_bnr_6')
// (7, 6, 'neigh_op_top_6')
// (7, 7, 'local_g1_6')
// (7, 7, 'lutff_3/in_0')
// (7, 7, 'lutff_6/out')
// (7, 8, 'neigh_op_bot_6')
// (8, 6, 'neigh_op_tnl_6')
// (8, 7, 'neigh_op_lft_6')
// (8, 8, 'neigh_op_bnl_6')

reg n371 = 0;
// (6, 7, 'neigh_op_tnr_0')
// (6, 8, 'neigh_op_rgt_0')
// (6, 9, 'neigh_op_bnr_0')
// (7, 7, 'neigh_op_top_0')
// (7, 8, 'local_g3_0')
// (7, 8, 'lutff_0/out')
// (7, 8, 'lutff_6/in_1')
// (7, 9, 'local_g0_0')
// (7, 9, 'lutff_0/in_2')
// (7, 9, 'neigh_op_bot_0')
// (8, 7, 'neigh_op_tnl_0')
// (8, 8, 'neigh_op_lft_0')
// (8, 9, 'neigh_op_bnl_0')

reg n372 = 0;
// (6, 7, 'neigh_op_tnr_1')
// (6, 8, 'neigh_op_rgt_1')
// (6, 9, 'neigh_op_bnr_1')
// (7, 7, 'neigh_op_top_1')
// (7, 8, 'local_g0_1')
// (7, 8, 'lutff_1/out')
// (7, 8, 'lutff_4/in_1')
// (7, 9, 'neigh_op_bot_1')
// (8, 7, 'neigh_op_tnl_1')
// (8, 8, 'neigh_op_lft_1')
// (8, 9, 'neigh_op_bnl_1')

reg n373 = 0;
// (6, 7, 'neigh_op_tnr_2')
// (6, 8, 'neigh_op_rgt_2')
// (6, 9, 'neigh_op_bnr_2')
// (7, 7, 'neigh_op_top_2')
// (7, 8, 'local_g0_2')
// (7, 8, 'local_g1_2')
// (7, 8, 'lutff_1/in_2')
// (7, 8, 'lutff_2/out')
// (7, 8, 'lutff_5/in_1')
// (7, 9, 'neigh_op_bot_2')
// (8, 7, 'neigh_op_tnl_2')
// (8, 8, 'neigh_op_lft_2')
// (8, 9, 'neigh_op_bnl_2')

reg n374 = 0;
// (6, 7, 'neigh_op_tnr_4')
// (6, 8, 'neigh_op_rgt_4')
// (6, 9, 'neigh_op_bnr_4')
// (7, 7, 'neigh_op_top_4')
// (7, 8, 'lutff_4/out')
// (7, 9, 'local_g1_4')
// (7, 9, 'lutff_0/in_1')
// (7, 9, 'neigh_op_bot_4')
// (8, 7, 'neigh_op_tnl_4')
// (8, 8, 'neigh_op_lft_4')
// (8, 9, 'neigh_op_bnl_4')

reg n375 = 0;
// (6, 7, 'neigh_op_tnr_5')
// (6, 8, 'neigh_op_rgt_5')
// (6, 9, 'neigh_op_bnr_5')
// (7, 7, 'neigh_op_top_5')
// (7, 8, 'local_g0_5')
// (7, 8, 'local_g1_5')
// (7, 8, 'lutff_0/in_1')
// (7, 8, 'lutff_4/in_2')
// (7, 8, 'lutff_5/out')
// (7, 9, 'neigh_op_bot_5')
// (8, 7, 'neigh_op_tnl_5')
// (8, 8, 'neigh_op_lft_5')
// (8, 9, 'neigh_op_bnl_5')

reg n376 = 0;
// (6, 7, 'neigh_op_tnr_6')
// (6, 8, 'local_g2_6')
// (6, 8, 'lutff_6/in_0')
// (6, 8, 'neigh_op_rgt_6')
// (6, 9, 'neigh_op_bnr_6')
// (7, 7, 'neigh_op_top_6')
// (7, 8, 'local_g1_6')
// (7, 8, 'lutff_2/in_1')
// (7, 8, 'lutff_6/out')
// (7, 9, 'neigh_op_bot_6')
// (8, 7, 'neigh_op_tnl_6')
// (8, 8, 'neigh_op_lft_6')
// (8, 9, 'neigh_op_bnl_6')

reg n377 = 0;
// (6, 7, 'neigh_op_tnr_7')
// (6, 7, 'sp4_r_v_b_43')
// (6, 8, 'neigh_op_rgt_7')
// (6, 8, 'sp4_r_v_b_30')
// (6, 9, 'neigh_op_bnr_7')
// (6, 9, 'sp4_r_v_b_19')
// (6, 10, 'sp4_r_v_b_6')
// (7, 6, 'sp4_v_t_43')
// (7, 7, 'neigh_op_top_7')
// (7, 7, 'sp4_v_b_43')
// (7, 8, 'lutff_7/out')
// (7, 8, 'sp4_v_b_30')
// (7, 9, 'neigh_op_bot_7')
// (7, 9, 'sp4_v_b_19')
// (7, 10, 'local_g0_6')
// (7, 10, 'lutff_2/in_0')
// (7, 10, 'sp4_v_b_6')
// (8, 7, 'neigh_op_tnl_7')
// (8, 8, 'neigh_op_lft_7')
// (8, 9, 'neigh_op_bnl_7')

reg n378 = 0;
// (6, 7, 'sp4_r_v_b_39')
// (6, 7, 'sp4_r_v_b_45')
// (6, 8, 'local_g0_3')
// (6, 8, 'lutff_3/in_2')
// (6, 8, 'sp4_r_v_b_26')
// (6, 8, 'sp4_r_v_b_32')
// (6, 9, 'sp4_r_v_b_15')
// (6, 9, 'sp4_r_v_b_21')
// (6, 10, 'sp4_r_v_b_2')
// (6, 10, 'sp4_r_v_b_8')
// (7, 6, 'sp4_h_r_8')
// (7, 6, 'sp4_v_t_39')
// (7, 6, 'sp4_v_t_45')
// (7, 7, 'sp4_v_b_39')
// (7, 7, 'sp4_v_b_45')
// (7, 8, 'local_g3_2')
// (7, 8, 'lutff_7/in_2')
// (7, 8, 'sp4_v_b_26')
// (7, 8, 'sp4_v_b_32')
// (7, 9, 'sp4_v_b_15')
// (7, 9, 'sp4_v_b_21')
// (7, 10, 'sp4_v_b_2')
// (7, 10, 'sp4_v_b_8')
// (8, 5, 'neigh_op_tnr_0')
// (8, 6, 'local_g3_0')
// (8, 6, 'lutff_5/in_0')
// (8, 6, 'neigh_op_rgt_0')
// (8, 6, 'sp4_h_r_21')
// (8, 7, 'neigh_op_bnr_0')
// (9, 5, 'neigh_op_top_0')
// (9, 6, 'lutff_0/out')
// (9, 6, 'sp4_h_r_32')
// (9, 7, 'local_g1_0')
// (9, 7, 'lutff_3/in_0')
// (9, 7, 'neigh_op_bot_0')
// (10, 5, 'neigh_op_tnl_0')
// (10, 6, 'neigh_op_lft_0')
// (10, 6, 'sp4_h_r_45')
// (10, 7, 'neigh_op_bnl_0')
// (11, 6, 'sp4_h_l_45')

wire n379;
// (6, 8, 'neigh_op_tnr_0')
// (6, 9, 'neigh_op_rgt_0')
// (6, 10, 'neigh_op_bnr_0')
// (7, 8, 'neigh_op_top_0')
// (7, 9, 'lutff_0/out')
// (7, 10, 'neigh_op_bot_0')
// (8, 8, 'neigh_op_tnl_0')
// (8, 9, 'local_g0_0')
// (8, 9, 'local_g1_0')
// (8, 9, 'lutff_0/in_1')
// (8, 9, 'lutff_3/in_1')
// (8, 9, 'neigh_op_lft_0')
// (8, 10, 'neigh_op_bnl_0')

reg n380 = 0;
// (6, 8, 'neigh_op_tnr_1')
// (6, 9, 'neigh_op_rgt_1')
// (6, 10, 'neigh_op_bnr_1')
// (7, 8, 'neigh_op_top_1')
// (7, 9, 'local_g1_1')
// (7, 9, 'lutff_1/out')
// (7, 9, 'lutff_2/in_0')
// (7, 10, 'neigh_op_bot_1')
// (8, 8, 'neigh_op_tnl_1')
// (8, 9, 'neigh_op_lft_1')
// (8, 10, 'neigh_op_bnl_1')

reg n381 = 0;
// (6, 8, 'neigh_op_tnr_2')
// (6, 9, 'neigh_op_rgt_2')
// (6, 10, 'neigh_op_bnr_2')
// (7, 8, 'neigh_op_top_2')
// (7, 9, 'local_g1_2')
// (7, 9, 'lutff_2/out')
// (7, 9, 'lutff_3/in_0')
// (7, 10, 'neigh_op_bot_2')
// (8, 8, 'neigh_op_tnl_2')
// (8, 9, 'neigh_op_lft_2')
// (8, 10, 'neigh_op_bnl_2')

reg n382 = 0;
// (6, 8, 'neigh_op_tnr_3')
// (6, 9, 'neigh_op_rgt_3')
// (6, 10, 'neigh_op_bnr_3')
// (7, 8, 'neigh_op_top_3')
// (7, 9, 'local_g1_3')
// (7, 9, 'lutff_3/out')
// (7, 9, 'lutff_4/in_0')
// (7, 10, 'neigh_op_bot_3')
// (8, 8, 'neigh_op_tnl_3')
// (8, 9, 'neigh_op_lft_3')
// (8, 10, 'neigh_op_bnl_3')

reg n383 = 0;
// (6, 8, 'neigh_op_tnr_7')
// (6, 9, 'neigh_op_rgt_7')
// (6, 10, 'neigh_op_bnr_7')
// (7, 8, 'neigh_op_top_7')
// (7, 9, 'local_g0_7')
// (7, 9, 'lutff_5/in_0')
// (7, 9, 'lutff_7/out')
// (7, 10, 'neigh_op_bot_7')
// (8, 8, 'neigh_op_tnl_7')
// (8, 9, 'neigh_op_lft_7')
// (8, 10, 'neigh_op_bnl_7')

wire n384;
// (6, 9, 'neigh_op_tnr_0')
// (6, 10, 'neigh_op_rgt_0')
// (6, 11, 'neigh_op_bnr_0')
// (7, 0, 'span12_vert_19')
// (7, 1, 'sp12_v_b_19')
// (7, 2, 'sp12_v_b_16')
// (7, 3, 'sp12_v_b_15')
// (7, 4, 'sp12_v_b_12')
// (7, 5, 'sp12_v_b_11')
// (7, 6, 'local_g3_0')
// (7, 6, 'lutff_0/in_3')
// (7, 6, 'sp12_v_b_8')
// (7, 7, 'sp12_v_b_7')
// (7, 8, 'sp12_v_b_4')
// (7, 9, 'neigh_op_top_0')
// (7, 9, 'sp12_v_b_3')
// (7, 10, 'lutff_0/out')
// (7, 10, 'sp12_v_b_0')
// (7, 11, 'neigh_op_bot_0')
// (8, 9, 'neigh_op_tnl_0')
// (8, 10, 'neigh_op_lft_0')
// (8, 11, 'neigh_op_bnl_0')

reg n385 = 0;
// (6, 9, 'neigh_op_tnr_5')
// (6, 9, 'sp4_r_v_b_39')
// (6, 10, 'neigh_op_rgt_5')
// (6, 10, 'sp4_r_v_b_26')
// (6, 11, 'neigh_op_bnr_5')
// (6, 11, 'sp4_r_v_b_15')
// (6, 12, 'sp4_r_v_b_2')
// (7, 8, 'sp4_h_r_2')
// (7, 8, 'sp4_v_t_39')
// (7, 9, 'neigh_op_top_5')
// (7, 9, 'sp4_v_b_39')
// (7, 10, 'local_g1_5')
// (7, 10, 'lutff_0/in_2')
// (7, 10, 'lutff_5/out')
// (7, 10, 'sp4_v_b_26')
// (7, 11, 'neigh_op_bot_5')
// (7, 11, 'sp4_v_b_15')
// (7, 12, 'local_g0_2')
// (7, 12, 'lutff_2/in_0')
// (7, 12, 'lutff_4/in_2')
// (7, 12, 'sp4_v_b_2')
// (8, 8, 'local_g0_7')
// (8, 8, 'lutff_3/in_0')
// (8, 8, 'sp4_h_r_15')
// (8, 9, 'neigh_op_tnl_5')
// (8, 10, 'neigh_op_lft_5')
// (8, 11, 'neigh_op_bnl_5')
// (9, 8, 'sp4_h_r_26')
// (10, 8, 'sp4_h_r_39')
// (11, 8, 'sp4_h_l_39')

reg n386 = 0;
// (6, 9, 'neigh_op_tnr_7')
// (6, 10, 'neigh_op_rgt_7')
// (6, 11, 'neigh_op_bnr_7')
// (7, 8, 'sp4_r_v_b_39')
// (7, 9, 'neigh_op_top_7')
// (7, 9, 'sp4_r_v_b_26')
// (7, 10, 'lutff_7/out')
// (7, 10, 'sp4_r_v_b_15')
// (7, 11, 'neigh_op_bot_7')
// (7, 11, 'sp4_r_v_b_2')
// (8, 7, 'sp4_v_t_39')
// (8, 8, 'sp4_v_b_39')
// (8, 9, 'neigh_op_tnl_7')
// (8, 9, 'sp4_v_b_26')
// (8, 10, 'neigh_op_lft_7')
// (8, 10, 'sp4_v_b_15')
// (8, 11, 'neigh_op_bnl_7')
// (8, 11, 'sp4_h_r_8')
// (8, 11, 'sp4_v_b_2')
// (9, 11, 'local_g1_5')
// (9, 11, 'lutff_0/in_2')
// (9, 11, 'sp4_h_r_21')
// (10, 11, 'sp4_h_r_32')
// (11, 11, 'sp4_h_r_45')
// (12, 11, 'sp4_h_l_45')

reg n387 = 0;
// (6, 9, 'sp12_h_r_1')
// (7, 9, 'sp12_h_r_2')
// (8, 8, 'neigh_op_tnr_7')
// (8, 9, 'neigh_op_rgt_7')
// (8, 9, 'sp12_h_r_5')
// (8, 10, 'neigh_op_bnr_7')
// (9, 8, 'neigh_op_top_7')
// (9, 9, 'lutff_7/out')
// (9, 9, 'sp12_h_r_6')
// (9, 10, 'neigh_op_bot_7')
// (10, 8, 'neigh_op_tnl_7')
// (10, 9, 'neigh_op_lft_7')
// (10, 9, 'sp12_h_r_9')
// (10, 10, 'neigh_op_bnl_7')
// (11, 9, 'local_g1_2')
// (11, 9, 'lutff_7/in_0')
// (11, 9, 'sp12_h_r_10')
// (12, 9, 'sp12_h_r_13')
// (13, 9, 'span12_horz_13')

reg n388 = 0;
// (6, 11, 'neigh_op_tnr_0')
// (6, 12, 'neigh_op_rgt_0')
// (6, 13, 'neigh_op_bnr_0')
// (7, 11, 'neigh_op_top_0')
// (7, 12, 'lutff_0/out')
// (7, 13, 'local_g1_0')
// (7, 13, 'lutff_7/in_0')
// (7, 13, 'neigh_op_bot_0')
// (8, 11, 'neigh_op_tnl_0')
// (8, 12, 'neigh_op_lft_0')
// (8, 13, 'neigh_op_bnl_0')

reg n389 = 0;
// (6, 11, 'neigh_op_tnr_1')
// (6, 12, 'neigh_op_rgt_1')
// (6, 13, 'neigh_op_bnr_1')
// (7, 11, 'neigh_op_top_1')
// (7, 12, 'local_g0_1')
// (7, 12, 'lutff_1/out')
// (7, 12, 'lutff_7/in_0')
// (7, 13, 'neigh_op_bot_1')
// (8, 11, 'neigh_op_tnl_1')
// (8, 12, 'neigh_op_lft_1')
// (8, 13, 'neigh_op_bnl_1')

reg n390 = 0;
// (6, 11, 'neigh_op_tnr_2')
// (6, 12, 'neigh_op_rgt_2')
// (6, 13, 'neigh_op_bnr_2')
// (7, 11, 'neigh_op_top_2')
// (7, 12, 'local_g1_2')
// (7, 12, 'lutff_1/in_0')
// (7, 12, 'lutff_2/out')
// (7, 13, 'neigh_op_bot_2')
// (8, 11, 'neigh_op_tnl_2')
// (8, 12, 'neigh_op_lft_2')
// (8, 13, 'neigh_op_bnl_2')

reg n391 = 0;
// (6, 11, 'neigh_op_tnr_4')
// (6, 12, 'neigh_op_rgt_4')
// (6, 13, 'neigh_op_bnr_4')
// (7, 11, 'neigh_op_top_4')
// (7, 12, 'local_g0_4')
// (7, 12, 'lutff_4/out')
// (7, 12, 'lutff_6/in_0')
// (7, 13, 'neigh_op_bot_4')
// (8, 11, 'neigh_op_tnl_4')
// (8, 12, 'neigh_op_lft_4')
// (8, 13, 'neigh_op_bnl_4')

reg n392 = 0;
// (6, 11, 'neigh_op_tnr_5')
// (6, 12, 'local_g3_5')
// (6, 12, 'lutff_2/in_0')
// (6, 12, 'neigh_op_rgt_5')
// (6, 13, 'neigh_op_bnr_5')
// (7, 11, 'neigh_op_top_5')
// (7, 12, 'lutff_5/out')
// (7, 13, 'neigh_op_bot_5')
// (8, 11, 'neigh_op_tnl_5')
// (8, 12, 'neigh_op_lft_5')
// (8, 13, 'neigh_op_bnl_5')

reg n393 = 0;
// (6, 11, 'neigh_op_tnr_6')
// (6, 12, 'neigh_op_rgt_6')
// (6, 13, 'neigh_op_bnr_6')
// (7, 11, 'neigh_op_top_6')
// (7, 12, 'local_g0_6')
// (7, 12, 'lutff_0/in_0')
// (7, 12, 'lutff_6/out')
// (7, 13, 'neigh_op_bot_6')
// (8, 11, 'neigh_op_tnl_6')
// (8, 12, 'neigh_op_lft_6')
// (8, 13, 'neigh_op_bnl_6')

reg n394 = 0;
// (6, 11, 'neigh_op_tnr_7')
// (6, 12, 'neigh_op_rgt_7')
// (6, 13, 'neigh_op_bnr_7')
// (7, 11, 'neigh_op_top_7')
// (7, 12, 'local_g2_7')
// (7, 12, 'lutff_5/in_0')
// (7, 12, 'lutff_7/out')
// (7, 13, 'neigh_op_bot_7')
// (8, 11, 'neigh_op_tnl_7')
// (8, 12, 'neigh_op_lft_7')
// (8, 13, 'neigh_op_bnl_7')

reg n395 = 0;
// (6, 11, 'sp4_h_r_7')
// (7, 11, 'local_g0_2')
// (7, 11, 'lutff_5/in_3')
// (7, 11, 'sp4_h_r_18')
// (8, 11, 'sp4_h_r_31')
// (9, 11, 'local_g3_2')
// (9, 11, 'lutff_0/in_1')
// (9, 11, 'sp4_h_r_42')
// (10, 10, 'neigh_op_tnr_3')
// (10, 11, 'neigh_op_rgt_3')
// (10, 11, 'sp4_h_l_42')
// (10, 11, 'sp4_h_r_11')
// (10, 12, 'neigh_op_bnr_3')
// (11, 10, 'neigh_op_top_3')
// (11, 11, 'lutff_3/out')
// (11, 11, 'sp4_h_r_22')
// (11, 12, 'neigh_op_bot_3')
// (12, 10, 'neigh_op_tnl_3')
// (12, 11, 'neigh_op_lft_3')
// (12, 11, 'sp4_h_r_35')
// (12, 12, 'neigh_op_bnl_3')
// (13, 11, 'span4_horz_35')

wire n396;
// (6, 12, 'neigh_op_tnr_0')
// (6, 13, 'neigh_op_rgt_0')
// (6, 14, 'neigh_op_bnr_0')
// (7, 12, 'neigh_op_top_0')
// (7, 13, 'local_g2_0')
// (7, 13, 'lutff_0/out')
// (7, 13, 'lutff_1/in_3')
// (7, 14, 'neigh_op_bot_0')
// (8, 12, 'neigh_op_tnl_0')
// (8, 13, 'neigh_op_lft_0')
// (8, 14, 'neigh_op_bnl_0')

wire n397;
// (6, 12, 'neigh_op_tnr_1')
// (6, 13, 'neigh_op_rgt_1')
// (6, 14, 'neigh_op_bnr_1')
// (7, 2, 'sp12_v_t_22')
// (7, 3, 'sp12_v_b_22')
// (7, 4, 'sp12_v_b_21')
// (7, 5, 'sp12_v_b_18')
// (7, 6, 'sp12_v_b_17')
// (7, 7, 'sp12_v_b_14')
// (7, 8, 'sp12_v_b_13')
// (7, 9, 'sp12_v_b_10')
// (7, 10, 'local_g2_1')
// (7, 10, 'lutff_0/in_3')
// (7, 10, 'sp12_v_b_9')
// (7, 11, 'sp12_v_b_6')
// (7, 12, 'neigh_op_top_1')
// (7, 12, 'sp12_v_b_5')
// (7, 13, 'lutff_1/out')
// (7, 13, 'sp12_v_b_2')
// (7, 14, 'neigh_op_bot_1')
// (7, 14, 'sp12_v_b_1')
// (8, 12, 'neigh_op_tnl_1')
// (8, 13, 'neigh_op_lft_1')
// (8, 14, 'neigh_op_bnl_1')

reg n398 = 0;
// (6, 12, 'neigh_op_tnr_2')
// (6, 13, 'neigh_op_rgt_2')
// (6, 14, 'neigh_op_bnr_2')
// (7, 12, 'neigh_op_top_2')
// (7, 13, 'local_g0_2')
// (7, 13, 'lutff_0/in_0')
// (7, 13, 'lutff_2/out')
// (7, 13, 'sp4_r_v_b_37')
// (7, 14, 'local_g0_0')
// (7, 14, 'lutff_5/in_1')
// (7, 14, 'neigh_op_bot_2')
// (7, 14, 'sp4_r_v_b_24')
// (7, 15, 'sp4_r_v_b_13')
// (7, 16, 'sp4_r_v_b_0')
// (8, 12, 'neigh_op_tnl_2')
// (8, 12, 'sp4_v_t_37')
// (8, 13, 'neigh_op_lft_2')
// (8, 13, 'sp4_v_b_37')
// (8, 14, 'neigh_op_bnl_2')
// (8, 14, 'sp4_v_b_24')
// (8, 15, 'sp4_v_b_13')
// (8, 16, 'sp4_v_b_0')

reg n399 = 0;
// (6, 12, 'neigh_op_tnr_4')
// (6, 13, 'neigh_op_rgt_4')
// (6, 14, 'neigh_op_bnr_4')
// (7, 12, 'neigh_op_top_4')
// (7, 13, 'local_g3_4')
// (7, 13, 'lutff_4/out')
// (7, 13, 'lutff_5/in_0')
// (7, 14, 'neigh_op_bot_4')
// (8, 12, 'neigh_op_tnl_4')
// (8, 13, 'neigh_op_lft_4')
// (8, 14, 'neigh_op_bnl_4')

reg n400 = 0;
// (6, 12, 'neigh_op_tnr_5')
// (6, 13, 'neigh_op_rgt_5')
// (6, 14, 'neigh_op_bnr_5')
// (7, 12, 'neigh_op_top_5')
// (7, 13, 'local_g3_5')
// (7, 13, 'lutff_2/in_0')
// (7, 13, 'lutff_5/out')
// (7, 14, 'neigh_op_bot_5')
// (8, 12, 'neigh_op_tnl_5')
// (8, 13, 'neigh_op_lft_5')
// (8, 14, 'neigh_op_bnl_5')

reg n401 = 0;
// (6, 12, 'neigh_op_tnr_6')
// (6, 13, 'neigh_op_rgt_6')
// (6, 14, 'neigh_op_bnr_6')
// (7, 12, 'neigh_op_top_6')
// (7, 13, 'local_g0_6')
// (7, 13, 'lutff_4/in_0')
// (7, 13, 'lutff_6/out')
// (7, 14, 'neigh_op_bot_6')
// (8, 12, 'neigh_op_tnl_6')
// (8, 13, 'neigh_op_lft_6')
// (8, 14, 'neigh_op_bnl_6')

reg n402 = 0;
// (6, 12, 'neigh_op_tnr_7')
// (6, 13, 'neigh_op_rgt_7')
// (6, 14, 'neigh_op_bnr_7')
// (7, 12, 'neigh_op_top_7')
// (7, 13, 'local_g2_7')
// (7, 13, 'lutff_0/in_1')
// (7, 13, 'lutff_6/in_1')
// (7, 13, 'lutff_7/out')
// (7, 14, 'neigh_op_bot_7')
// (8, 12, 'neigh_op_tnl_7')
// (8, 13, 'neigh_op_lft_7')
// (8, 14, 'neigh_op_bnl_7')

reg n403 = 0;
// (6, 13, 'neigh_op_tnr_2')
// (6, 14, 'neigh_op_rgt_2')
// (6, 15, 'neigh_op_bnr_2')
// (7, 13, 'neigh_op_top_2')
// (7, 14, 'local_g0_2')
// (7, 14, 'lutff_2/out')
// (7, 14, 'lutff_6/in_0')
// (7, 15, 'neigh_op_bot_2')
// (8, 13, 'neigh_op_tnl_2')
// (8, 14, 'neigh_op_lft_2')
// (8, 15, 'neigh_op_bnl_2')

reg n404 = 0;
// (6, 13, 'neigh_op_tnr_5')
// (6, 14, 'neigh_op_rgt_5')
// (6, 15, 'neigh_op_bnr_5')
// (7, 13, 'neigh_op_top_5')
// (7, 14, 'local_g1_5')
// (7, 14, 'lutff_2/in_0')
// (7, 14, 'lutff_5/out')
// (7, 15, 'neigh_op_bot_5')
// (8, 13, 'neigh_op_tnl_5')
// (8, 14, 'neigh_op_lft_5')
// (8, 15, 'neigh_op_bnl_5')

reg n405 = 0;
// (6, 13, 'neigh_op_tnr_6')
// (6, 14, 'neigh_op_rgt_6')
// (6, 15, 'neigh_op_bnr_6')
// (7, 13, 'neigh_op_top_6')
// (7, 14, 'local_g1_6')
// (7, 14, 'lutff_6/out')
// (7, 14, 'lutff_7/in_0')
// (7, 15, 'neigh_op_bot_6')
// (8, 13, 'neigh_op_tnl_6')
// (8, 14, 'neigh_op_lft_6')
// (8, 15, 'neigh_op_bnl_6')

reg n406 = 0;
// (6, 13, 'neigh_op_tnr_7')
// (6, 14, 'neigh_op_rgt_7')
// (6, 15, 'neigh_op_bnr_7')
// (7, 9, 'sp12_v_t_22')
// (7, 10, 'sp12_v_b_22')
// (7, 11, 'sp12_v_b_21')
// (7, 12, 'local_g2_2')
// (7, 12, 'lutff_4/in_0')
// (7, 12, 'sp12_v_b_18')
// (7, 13, 'local_g0_7')
// (7, 13, 'local_g1_7')
// (7, 13, 'lutff_1/in_0')
// (7, 13, 'lutff_6/in_0')
// (7, 13, 'neigh_op_top_7')
// (7, 13, 'sp12_v_b_17')
// (7, 14, 'local_g0_7')
// (7, 14, 'lutff_5/in_0')
// (7, 14, 'lutff_7/out')
// (7, 14, 'sp12_v_b_14')
// (7, 15, 'neigh_op_bot_7')
// (7, 15, 'sp12_v_b_13')
// (7, 16, 'sp12_v_b_10')
// (7, 17, 'span12_vert_9')
// (8, 13, 'neigh_op_tnl_7')
// (8, 14, 'neigh_op_lft_7')
// (8, 15, 'neigh_op_bnl_7')

wire n407;
// (7, 1, 'local_g3_5')
// (7, 1, 'lutff_1/in_3')
// (7, 1, 'lutff_3/in_3')
// (7, 1, 'neigh_op_tnr_5')
// (7, 2, 'neigh_op_rgt_5')
// (7, 3, 'neigh_op_bnr_5')
// (8, 1, 'neigh_op_top_5')
// (8, 2, 'local_g1_5')
// (8, 2, 'lutff_0/in_0')
// (8, 2, 'lutff_5/out')
// (8, 3, 'neigh_op_bot_5')
// (9, 1, 'neigh_op_tnl_5')
// (9, 2, 'neigh_op_lft_5')
// (9, 3, 'neigh_op_bnl_5')

wire n408;
// (7, 1, 'neigh_op_tnr_0')
// (7, 2, 'local_g2_0')
// (7, 2, 'lutff_0/in_2')
// (7, 2, 'lutff_5/in_3')
// (7, 2, 'neigh_op_rgt_0')
// (7, 3, 'neigh_op_bnr_0')
// (8, 1, 'neigh_op_top_0')
// (8, 2, 'lutff_0/out')
// (8, 3, 'neigh_op_bot_0')
// (9, 1, 'neigh_op_tnl_0')
// (9, 2, 'neigh_op_lft_0')
// (9, 3, 'neigh_op_bnl_0')

wire n409;
// (7, 1, 'neigh_op_tnr_1')
// (7, 2, 'neigh_op_rgt_1')
// (7, 3, 'neigh_op_bnr_1')
// (8, 1, 'neigh_op_top_1')
// (8, 2, 'local_g2_1')
// (8, 2, 'lutff_1/out')
// (8, 2, 'lutff_2/in_3')
// (8, 3, 'neigh_op_bot_1')
// (9, 1, 'neigh_op_tnl_1')
// (9, 2, 'neigh_op_lft_1')
// (9, 3, 'neigh_op_bnl_1')

wire n410;
// (7, 1, 'neigh_op_tnr_3')
// (7, 2, 'neigh_op_rgt_3')
// (7, 3, 'neigh_op_bnr_3')
// (8, 1, 'neigh_op_top_3')
// (8, 2, 'local_g0_3')
// (8, 2, 'lutff_0/in_3')
// (8, 2, 'lutff_3/out')
// (8, 3, 'neigh_op_bot_3')
// (9, 1, 'neigh_op_tnl_3')
// (9, 2, 'neigh_op_lft_3')
// (9, 3, 'neigh_op_bnl_3')

wire n411;
// (7, 1, 'neigh_op_tnr_4')
// (7, 2, 'local_g3_4')
// (7, 2, 'lutff_0/in_3')
// (7, 2, 'lutff_4/in_3')
// (7, 2, 'neigh_op_rgt_4')
// (7, 3, 'neigh_op_bnr_4')
// (8, 1, 'neigh_op_top_4')
// (8, 2, 'lutff_4/out')
// (8, 3, 'neigh_op_bot_4')
// (9, 1, 'neigh_op_tnl_4')
// (9, 2, 'neigh_op_lft_4')
// (9, 3, 'neigh_op_bnl_4')

wire n412;
// (7, 1, 'neigh_op_tnr_7')
// (7, 2, 'neigh_op_rgt_7')
// (7, 3, 'neigh_op_bnr_7')
// (8, 1, 'neigh_op_top_7')
// (8, 2, 'local_g0_7')
// (8, 2, 'lutff_4/in_3')
// (8, 2, 'lutff_7/out')
// (8, 3, 'neigh_op_bot_7')
// (9, 1, 'neigh_op_tnl_7')
// (9, 2, 'neigh_op_lft_7')
// (9, 3, 'neigh_op_bnl_7')

wire n413;
// (7, 1, 'sp4_r_v_b_15')
// (7, 2, 'local_g1_2')
// (7, 2, 'local_g2_6')
// (7, 2, 'lutff_1/in_3')
// (7, 2, 'lutff_7/in_2')
// (7, 2, 'sp4_r_v_b_2')
// (7, 2, 'sp4_r_v_b_38')
// (7, 3, 'local_g3_7')
// (7, 3, 'lutff_4/in_2')
// (7, 3, 'lutff_6/in_2')
// (7, 3, 'neigh_op_tnr_7')
// (7, 3, 'sp4_r_v_b_27')
// (7, 3, 'sp4_r_v_b_43')
// (7, 4, 'neigh_op_rgt_7')
// (7, 4, 'sp4_r_v_b_14')
// (7, 4, 'sp4_r_v_b_30')
// (7, 5, 'neigh_op_bnr_7')
// (7, 5, 'sp4_r_v_b_19')
// (7, 5, 'sp4_r_v_b_3')
// (7, 6, 'sp4_r_v_b_6')
// (8, 0, 'span4_vert_15')
// (8, 1, 'sp4_v_b_15')
// (8, 1, 'sp4_v_t_38')
// (8, 2, 'local_g2_6')
// (8, 2, 'lutff_3/in_1')
// (8, 2, 'sp4_v_b_2')
// (8, 2, 'sp4_v_b_38')
// (8, 2, 'sp4_v_t_43')
// (8, 3, 'neigh_op_top_7')
// (8, 3, 'sp4_v_b_27')
// (8, 3, 'sp4_v_b_43')
// (8, 4, 'lutff_7/out')
// (8, 4, 'sp4_v_b_14')
// (8, 4, 'sp4_v_b_30')
// (8, 5, 'neigh_op_bot_7')
// (8, 5, 'sp4_v_b_19')
// (8, 5, 'sp4_v_b_3')
// (8, 6, 'sp4_v_b_6')
// (9, 3, 'neigh_op_tnl_7')
// (9, 4, 'neigh_op_lft_7')
// (9, 5, 'neigh_op_bnl_7')

wire n414;
// (7, 1, 'sp4_r_v_b_37')
// (7, 2, 'sp4_r_v_b_24')
// (7, 3, 'neigh_op_tnr_0')
// (7, 3, 'sp4_r_v_b_13')
// (7, 4, 'neigh_op_rgt_0')
// (7, 4, 'sp4_r_v_b_0')
// (7, 5, 'neigh_op_bnr_0')
// (8, 0, 'span4_vert_37')
// (8, 1, 'sp4_r_v_b_36')
// (8, 1, 'sp4_v_b_37')
// (8, 2, 'local_g0_1')
// (8, 2, 'local_g3_0')
// (8, 2, 'lutff_3/in_2')
// (8, 2, 'lutff_6/in_3')
// (8, 2, 'sp4_r_v_b_25')
// (8, 2, 'sp4_v_b_24')
// (8, 3, 'local_g1_0')
// (8, 3, 'lutff_6/in_3')
// (8, 3, 'neigh_op_top_0')
// (8, 3, 'sp4_r_v_b_12')
// (8, 3, 'sp4_v_b_13')
// (8, 4, 'lutff_0/out')
// (8, 4, 'sp4_r_v_b_1')
// (8, 4, 'sp4_v_b_0')
// (8, 5, 'neigh_op_bot_0')
// (9, 0, 'span4_vert_36')
// (9, 1, 'sp4_v_b_36')
// (9, 2, 'sp4_v_b_25')
// (9, 3, 'neigh_op_tnl_0')
// (9, 3, 'sp4_v_b_12')
// (9, 4, 'neigh_op_lft_0')
// (9, 4, 'sp4_v_b_1')
// (9, 5, 'neigh_op_bnl_0')

wire n415;
// (7, 1, 'sp4_r_v_b_40')
// (7, 2, 'local_g1_5')
// (7, 2, 'lutff_2/in_2')
// (7, 2, 'lutff_3/in_1')
// (7, 2, 'neigh_op_tnr_0')
// (7, 2, 'sp4_r_v_b_29')
// (7, 3, 'neigh_op_rgt_0')
// (7, 3, 'sp4_r_v_b_16')
// (7, 4, 'neigh_op_bnr_0')
// (7, 4, 'sp4_r_v_b_5')
// (8, 0, 'span4_vert_40')
// (8, 1, 'sp4_v_b_40')
// (8, 2, 'local_g1_0')
// (8, 2, 'lutff_5/in_2')
// (8, 2, 'neigh_op_top_0')
// (8, 2, 'sp4_v_b_29')
// (8, 3, 'lutff_0/out')
// (8, 3, 'sp4_v_b_16')
// (8, 4, 'neigh_op_bot_0')
// (8, 4, 'sp4_v_b_5')
// (9, 2, 'neigh_op_tnl_0')
// (9, 3, 'neigh_op_lft_0')
// (9, 4, 'neigh_op_bnl_0')

wire n416;
// (7, 1, 'sp4_r_v_b_41')
// (7, 2, 'sp4_r_v_b_28')
// (7, 3, 'neigh_op_tnr_2')
// (7, 3, 'sp4_r_v_b_17')
// (7, 4, 'neigh_op_rgt_2')
// (7, 4, 'sp4_r_v_b_4')
// (7, 5, 'neigh_op_bnr_2')
// (8, 0, 'span4_vert_41')
// (8, 1, 'sp4_r_v_b_40')
// (8, 1, 'sp4_v_b_41')
// (8, 2, 'local_g0_5')
// (8, 2, 'local_g2_4')
// (8, 2, 'lutff_1/in_2')
// (8, 2, 'lutff_7/in_1')
// (8, 2, 'sp4_r_v_b_29')
// (8, 2, 'sp4_v_b_28')
// (8, 3, 'local_g1_1')
// (8, 3, 'lutff_5/in_3')
// (8, 3, 'neigh_op_top_2')
// (8, 3, 'sp4_r_v_b_16')
// (8, 3, 'sp4_v_b_17')
// (8, 4, 'local_g1_2')
// (8, 4, 'lutff_2/out')
// (8, 4, 'lutff_7/in_2')
// (8, 4, 'sp4_r_v_b_5')
// (8, 4, 'sp4_v_b_4')
// (8, 5, 'neigh_op_bot_2')
// (9, 0, 'span4_vert_40')
// (9, 1, 'sp4_v_b_40')
// (9, 2, 'sp4_v_b_29')
// (9, 3, 'neigh_op_tnl_2')
// (9, 3, 'sp4_v_b_16')
// (9, 4, 'neigh_op_lft_2')
// (9, 4, 'sp4_v_b_5')
// (9, 5, 'neigh_op_bnl_2')

wire n417;
// (7, 2, 'local_g2_4')
// (7, 2, 'lutff_1/in_1')
// (7, 2, 'lutff_7/in_3')
// (7, 2, 'neigh_op_tnr_4')
// (7, 3, 'local_g2_4')
// (7, 3, 'local_g3_4')
// (7, 3, 'lutff_3/in_1')
// (7, 3, 'lutff_5/in_2')
// (7, 3, 'neigh_op_rgt_4')
// (7, 4, 'neigh_op_bnr_4')
// (8, 2, 'local_g0_4')
// (8, 2, 'local_g1_4')
// (8, 2, 'lutff_3/in_0')
// (8, 2, 'lutff_6/in_2')
// (8, 2, 'neigh_op_top_4')
// (8, 3, 'local_g0_4')
// (8, 3, 'lutff_4/out')
// (8, 3, 'lutff_6/in_2')
// (8, 4, 'neigh_op_bot_4')
// (9, 2, 'neigh_op_tnl_4')
// (9, 3, 'neigh_op_lft_4')
// (9, 4, 'neigh_op_bnl_4')

wire n418;
// (7, 2, 'local_g3_6')
// (7, 2, 'lutff_1/in_2')
// (7, 2, 'lutff_2/in_1')
// (7, 2, 'neigh_op_tnr_6')
// (7, 3, 'local_g3_6')
// (7, 3, 'lutff_4/in_3')
// (7, 3, 'lutff_6/in_3')
// (7, 3, 'neigh_op_rgt_6')
// (7, 4, 'neigh_op_bnr_6')
// (8, 2, 'local_g1_6')
// (8, 2, 'lutff_2/in_1')
// (8, 2, 'neigh_op_top_6')
// (8, 3, 'lutff_6/out')
// (8, 4, 'neigh_op_bot_6')
// (9, 2, 'neigh_op_tnl_6')
// (9, 3, 'neigh_op_lft_6')
// (9, 4, 'neigh_op_bnl_6')

reg n419 = 0;
// (7, 2, 'sp4_r_v_b_36')
// (7, 3, 'sp4_r_v_b_25')
// (7, 4, 'sp4_r_v_b_12')
// (7, 5, 'sp4_r_v_b_1')
// (7, 6, 'sp4_h_r_6')
// (8, 0, 'span12_vert_6')
// (8, 1, 'sp12_v_b_6')
// (8, 1, 'sp4_v_t_36')
// (8, 2, 'sp12_v_b_5')
// (8, 2, 'sp4_v_b_36')
// (8, 3, 'sp12_v_b_2')
// (8, 3, 'sp4_v_b_25')
// (8, 4, 'sp12_h_r_1')
// (8, 4, 'sp12_v_b_1')
// (8, 4, 'sp12_v_t_22')
// (8, 4, 'sp4_v_b_12')
// (8, 5, 'local_g0_1')
// (8, 5, 'local_g2_6')
// (8, 5, 'lutff_0/in_0')
// (8, 5, 'lutff_1/in_0')
// (8, 5, 'lutff_3/in_0')
// (8, 5, 'sp12_v_b_22')
// (8, 5, 'sp4_h_r_1')
// (8, 5, 'sp4_v_b_1')
// (8, 6, 'local_g0_3')
// (8, 6, 'local_g3_5')
// (8, 6, 'lutff_0/in_0')
// (8, 6, 'lutff_1/in_0')
// (8, 6, 'lutff_2/in_0')
// (8, 6, 'lutff_3/in_0')
// (8, 6, 'lutff_4/in_0')
// (8, 6, 'sp12_v_b_21')
// (8, 6, 'sp4_h_r_19')
// (8, 7, 'local_g2_2')
// (8, 7, 'local_g3_2')
// (8, 7, 'lutff_0/in_1')
// (8, 7, 'lutff_1/in_0')
// (8, 7, 'lutff_3/in_0')
// (8, 7, 'lutff_4/in_0')
// (8, 7, 'sp12_v_b_18')
// (8, 8, 'sp12_v_b_17')
// (8, 9, 'sp12_v_b_14')
// (8, 10, 'sp12_v_b_13')
// (8, 11, 'sp12_v_b_10')
// (8, 12, 'sp12_v_b_9')
// (8, 13, 'sp12_v_b_6')
// (8, 14, 'sp12_v_b_5')
// (8, 15, 'sp12_v_b_2')
// (8, 16, 'sp12_v_b_1')
// (9, 4, 'local_g1_2')
// (9, 4, 'lutff_1/in_0')
// (9, 4, 'lutff_2/in_3')
// (9, 4, 'sp12_h_r_2')
// (9, 5, 'local_g0_4')
// (9, 5, 'lutff_1/in_3')
// (9, 5, 'sp4_h_r_12')
// (9, 6, 'sp4_h_r_30')
// (10, 3, 'neigh_op_tnr_7')
// (10, 3, 'sp4_r_v_b_43')
// (10, 4, 'neigh_op_rgt_7')
// (10, 4, 'sp12_h_r_5')
// (10, 4, 'sp4_r_v_b_30')
// (10, 5, 'neigh_op_bnr_7')
// (10, 5, 'sp4_h_r_25')
// (10, 5, 'sp4_r_v_b_19')
// (10, 6, 'sp4_h_r_43')
// (10, 6, 'sp4_r_v_b_6')
// (10, 7, 'sp4_r_v_b_44')
// (10, 8, 'sp4_r_v_b_33')
// (10, 9, 'sp4_r_v_b_20')
// (10, 10, 'sp4_r_v_b_9')
// (11, 2, 'sp4_v_t_43')
// (11, 3, 'neigh_op_top_7')
// (11, 3, 'sp4_v_b_43')
// (11, 4, 'local_g2_7')
// (11, 4, 'lutff_5/in_2')
// (11, 4, 'lutff_7/out')
// (11, 4, 'sp12_h_r_6')
// (11, 4, 'sp4_v_b_30')
// (11, 5, 'neigh_op_bot_7')
// (11, 5, 'sp4_h_r_36')
// (11, 5, 'sp4_v_b_19')
// (11, 6, 'local_g0_6')
// (11, 6, 'lutff_2/in_0')
// (11, 6, 'lutff_4/in_0')
// (11, 6, 'sp4_h_l_43')
// (11, 6, 'sp4_v_b_6')
// (11, 6, 'sp4_v_t_44')
// (11, 7, 'sp4_v_b_44')
// (11, 8, 'local_g2_1')
// (11, 8, 'lutff_1/in_2')
// (11, 8, 'sp4_v_b_33')
// (11, 9, 'sp4_v_b_20')
// (11, 10, 'sp4_v_b_9')
// (12, 3, 'neigh_op_tnl_7')
// (12, 4, 'neigh_op_lft_7')
// (12, 4, 'sp12_h_r_9')
// (12, 5, 'neigh_op_bnl_7')
// (12, 5, 'sp4_h_l_36')
// (13, 4, 'span12_horz_9')

wire n420;
// (7, 2, 'sp4_r_v_b_41')
// (7, 3, 'sp4_r_v_b_28')
// (7, 4, 'neigh_op_tnr_2')
// (7, 4, 'sp4_r_v_b_17')
// (7, 5, 'neigh_op_rgt_2')
// (7, 5, 'sp4_r_v_b_4')
// (7, 6, 'neigh_op_bnr_2')
// (8, 1, 'sp4_v_t_41')
// (8, 2, 'sp4_v_b_41')
// (8, 3, 'local_g2_4')
// (8, 3, 'local_g3_4')
// (8, 3, 'lutff_4/in_3')
// (8, 3, 'lutff_7/in_3')
// (8, 3, 'sp4_r_v_b_45')
// (8, 3, 'sp4_v_b_28')
// (8, 4, 'local_g2_0')
// (8, 4, 'lutff_3/in_1')
// (8, 4, 'neigh_op_top_2')
// (8, 4, 'sp4_r_v_b_32')
// (8, 4, 'sp4_v_b_17')
// (8, 5, 'lutff_2/out')
// (8, 5, 'sp4_r_v_b_21')
// (8, 5, 'sp4_v_b_4')
// (8, 6, 'neigh_op_bot_2')
// (8, 6, 'sp4_r_v_b_8')
// (9, 2, 'sp4_v_t_45')
// (9, 3, 'sp4_v_b_45')
// (9, 4, 'neigh_op_tnl_2')
// (9, 4, 'sp4_v_b_32')
// (9, 5, 'neigh_op_lft_2')
// (9, 5, 'sp4_v_b_21')
// (9, 6, 'neigh_op_bnl_2')
// (9, 6, 'sp4_v_b_8')

wire n421;
// (7, 3, 'neigh_op_tnr_3')
// (7, 4, 'neigh_op_rgt_3')
// (7, 5, 'neigh_op_bnr_3')
// (8, 0, 'span12_vert_13')
// (8, 1, 'sp12_v_b_13')
// (8, 2, 'local_g2_2')
// (8, 2, 'lutff_3/in_3')
// (8, 2, 'lutff_5/in_3')
// (8, 2, 'sp12_v_b_10')
// (8, 3, 'local_g1_3')
// (8, 3, 'lutff_1/in_3')
// (8, 3, 'neigh_op_top_3')
// (8, 3, 'sp12_v_b_9')
// (8, 4, 'lutff_3/out')
// (8, 4, 'sp12_v_b_6')
// (8, 4, 'sp4_h_r_6')
// (8, 5, 'neigh_op_bot_3')
// (8, 5, 'sp12_v_b_5')
// (8, 6, 'sp12_v_b_2')
// (8, 7, 'sp12_v_b_1')
// (9, 3, 'neigh_op_tnl_3')
// (9, 4, 'neigh_op_lft_3')
// (9, 4, 'sp4_h_r_19')
// (9, 5, 'neigh_op_bnl_3')
// (10, 4, 'sp4_h_r_30')
// (11, 1, 'sp4_r_v_b_37')
// (11, 2, 'local_g1_0')
// (11, 2, 'lutff_7/in_2')
// (11, 2, 'sp4_r_v_b_24')
// (11, 3, 'sp4_r_v_b_13')
// (11, 4, 'sp4_h_r_43')
// (11, 4, 'sp4_r_v_b_0')
// (12, 0, 'span4_vert_37')
// (12, 1, 'sp4_v_b_37')
// (12, 2, 'sp4_v_b_24')
// (12, 3, 'sp4_v_b_13')
// (12, 4, 'sp4_h_l_43')
// (12, 4, 'sp4_v_b_0')

wire n422;
// (7, 3, 'neigh_op_tnr_4')
// (7, 4, 'neigh_op_rgt_4')
// (7, 5, 'neigh_op_bnr_4')
// (8, 3, 'neigh_op_top_4')
// (8, 4, 'local_g0_4')
// (8, 4, 'local_g1_4')
// (8, 4, 'lutff_0/in_3')
// (8, 4, 'lutff_3/in_2')
// (8, 4, 'lutff_4/out')
// (8, 4, 'lutff_6/in_2')
// (8, 5, 'neigh_op_bot_4')
// (9, 3, 'neigh_op_tnl_4')
// (9, 4, 'neigh_op_lft_4')
// (9, 5, 'neigh_op_bnl_4')

wire n423;
// (7, 3, 'neigh_op_tnr_5')
// (7, 4, 'neigh_op_rgt_5')
// (7, 5, 'neigh_op_bnr_5')
// (8, 3, 'neigh_op_top_5')
// (8, 4, 'local_g3_5')
// (8, 4, 'lutff_3/in_3')
// (8, 4, 'lutff_5/out')
// (8, 5, 'neigh_op_bot_5')
// (9, 3, 'neigh_op_tnl_5')
// (9, 4, 'neigh_op_lft_5')
// (9, 5, 'neigh_op_bnl_5')

wire n424;
// (7, 3, 'sp4_h_r_9')
// (7, 3, 'sp4_r_v_b_36')
// (7, 4, 'sp4_r_v_b_25')
// (7, 5, 'sp4_r_v_b_12')
// (7, 6, 'sp4_r_v_b_1')
// (8, 2, 'sp4_v_t_36')
// (8, 3, 'local_g1_4')
// (8, 3, 'lutff_3/in_2')
// (8, 3, 'sp4_h_r_20')
// (8, 3, 'sp4_v_b_36')
// (8, 4, 'local_g3_1')
// (8, 4, 'lutff_4/in_0')
// (8, 4, 'sp4_v_b_25')
// (8, 5, 'local_g1_4')
// (8, 5, 'lutff_6/in_1')
// (8, 5, 'sp4_v_b_12')
// (8, 6, 'sp4_h_r_1')
// (8, 6, 'sp4_v_b_1')
// (9, 3, 'sp4_h_r_33')
// (9, 6, 'sp4_h_r_12')
// (10, 3, 'sp4_h_r_44')
// (10, 4, 'sp4_r_v_b_44')
// (10, 5, 'neigh_op_tnr_2')
// (10, 5, 'sp4_r_v_b_33')
// (10, 6, 'neigh_op_rgt_2')
// (10, 6, 'sp4_h_r_25')
// (10, 6, 'sp4_r_v_b_20')
// (10, 7, 'neigh_op_bnr_2')
// (10, 7, 'sp4_r_v_b_9')
// (11, 3, 'sp4_h_l_44')
// (11, 3, 'sp4_v_t_44')
// (11, 4, 'sp4_v_b_44')
// (11, 5, 'neigh_op_top_2')
// (11, 5, 'sp4_v_b_33')
// (11, 6, 'lutff_2/out')
// (11, 6, 'sp4_h_r_36')
// (11, 6, 'sp4_v_b_20')
// (11, 7, 'neigh_op_bot_2')
// (11, 7, 'sp4_v_b_9')
// (12, 5, 'neigh_op_tnl_2')
// (12, 6, 'neigh_op_lft_2')
// (12, 6, 'sp4_h_l_36')
// (12, 7, 'neigh_op_bnl_2')

reg n425 = 0;
// (7, 3, 'sp4_r_v_b_45')
// (7, 4, 'local_g0_3')
// (7, 4, 'lutff_0/in_3')
// (7, 4, 'sp4_r_v_b_32')
// (7, 5, 'sp4_r_v_b_21')
// (7, 6, 'sp4_r_v_b_8')
// (8, 2, 'sp4_v_t_45')
// (8, 3, 'sp4_v_b_45')
// (8, 4, 'sp4_v_b_32')
// (8, 5, 'sp4_v_b_21')
// (8, 6, 'sp4_h_r_8')
// (8, 6, 'sp4_v_b_8')
// (9, 6, 'sp4_h_r_21')
// (10, 6, 'sp4_h_r_32')
// (10, 8, 'neigh_op_tnr_2')
// (10, 9, 'neigh_op_rgt_2')
// (10, 10, 'neigh_op_bnr_2')
// (11, 6, 'sp4_h_r_45')
// (11, 7, 'sp4_r_v_b_45')
// (11, 8, 'neigh_op_top_2')
// (11, 8, 'sp4_r_v_b_32')
// (11, 9, 'lutff_2/out')
// (11, 9, 'sp4_r_v_b_21')
// (11, 10, 'local_g0_2')
// (11, 10, 'lutff_5/in_1')
// (11, 10, 'neigh_op_bot_2')
// (11, 10, 'sp4_r_v_b_8')
// (12, 6, 'sp4_h_l_45')
// (12, 6, 'sp4_v_t_45')
// (12, 7, 'sp4_v_b_45')
// (12, 8, 'neigh_op_tnl_2')
// (12, 8, 'sp4_v_b_32')
// (12, 9, 'neigh_op_lft_2')
// (12, 9, 'sp4_v_b_21')
// (12, 10, 'neigh_op_bnl_2')
// (12, 10, 'sp4_v_b_8')

wire n426;
// (7, 3, 'sp4_r_v_b_46')
// (7, 4, 'neigh_op_tnr_3')
// (7, 4, 'sp4_r_v_b_35')
// (7, 5, 'neigh_op_rgt_3')
// (7, 5, 'sp4_r_v_b_22')
// (7, 6, 'neigh_op_bnr_3')
// (7, 6, 'sp4_r_v_b_11')
// (8, 2, 'sp4_v_t_46')
// (8, 3, 'sp4_v_b_46')
// (8, 4, 'local_g2_3')
// (8, 4, 'local_g3_3')
// (8, 4, 'lutff_2/in_3')
// (8, 4, 'lutff_4/in_2')
// (8, 4, 'neigh_op_top_3')
// (8, 4, 'sp4_v_b_35')
// (8, 5, 'lutff_3/out')
// (8, 5, 'sp4_v_b_22')
// (8, 6, 'neigh_op_bot_3')
// (8, 6, 'sp4_v_b_11')
// (9, 4, 'neigh_op_tnl_3')
// (9, 5, 'neigh_op_lft_3')
// (9, 6, 'neigh_op_bnl_3')

wire n427;
// (7, 3, 'sp4_r_v_b_47')
// (7, 4, 'sp4_r_v_b_34')
// (7, 5, 'sp4_r_v_b_23')
// (7, 6, 'sp4_r_v_b_10')
// (8, 2, 'sp4_v_t_47')
// (8, 3, 'local_g3_7')
// (8, 3, 'lutff_3/in_3')
// (8, 3, 'sp4_v_b_47')
// (8, 4, 'local_g3_2')
// (8, 4, 'lutff_4/in_3')
// (8, 4, 'sp4_v_b_34')
// (8, 5, 'local_g1_7')
// (8, 5, 'lutff_6/in_2')
// (8, 5, 'sp4_v_b_23')
// (8, 6, 'sp4_h_r_5')
// (8, 6, 'sp4_v_b_10')
// (9, 6, 'sp4_h_r_16')
// (10, 5, 'neigh_op_tnr_4')
// (10, 6, 'neigh_op_rgt_4')
// (10, 6, 'sp4_h_r_29')
// (10, 7, 'neigh_op_bnr_4')
// (11, 5, 'neigh_op_top_4')
// (11, 6, 'lutff_4/out')
// (11, 6, 'sp4_h_r_40')
// (11, 7, 'neigh_op_bot_4')
// (12, 5, 'neigh_op_tnl_4')
// (12, 6, 'neigh_op_lft_4')
// (12, 6, 'sp4_h_l_40')
// (12, 7, 'neigh_op_bnl_4')

wire n428;
// (7, 4, 'neigh_op_tnr_0')
// (7, 5, 'neigh_op_rgt_0')
// (7, 6, 'neigh_op_bnr_0')
// (8, 2, 'sp4_r_v_b_36')
// (8, 3, 'sp4_r_v_b_25')
// (8, 4, 'local_g2_4')
// (8, 4, 'lutff_1/in_3')
// (8, 4, 'lutff_5/in_3')
// (8, 4, 'neigh_op_top_0')
// (8, 4, 'sp4_r_v_b_12')
// (8, 5, 'lutff_0/out')
// (8, 5, 'sp4_r_v_b_1')
// (8, 6, 'neigh_op_bot_0')
// (9, 1, 'sp4_v_t_36')
// (9, 2, 'sp4_v_b_36')
// (9, 3, 'sp4_v_b_25')
// (9, 4, 'neigh_op_tnl_0')
// (9, 4, 'sp4_v_b_12')
// (9, 5, 'neigh_op_lft_0')
// (9, 5, 'sp4_v_b_1')
// (9, 6, 'neigh_op_bnl_0')

wire n429;
// (7, 4, 'neigh_op_tnr_1')
// (7, 5, 'neigh_op_rgt_1')
// (7, 6, 'neigh_op_bnr_1')
// (8, 4, 'neigh_op_top_1')
// (8, 5, 'local_g1_1')
// (8, 5, 'lutff_1/out')
// (8, 5, 'lutff_2/in_0')
// (8, 5, 'lutff_4/in_2')
// (8, 6, 'neigh_op_bot_1')
// (9, 4, 'neigh_op_tnl_1')
// (9, 5, 'neigh_op_lft_1')
// (9, 6, 'neigh_op_bnl_1')

wire n430;
// (7, 4, 'neigh_op_tnr_4')
// (7, 5, 'neigh_op_rgt_4')
// (7, 6, 'neigh_op_bnr_4')
// (8, 2, 'sp4_r_v_b_44')
// (8, 3, 'local_g0_2')
// (8, 3, 'local_g2_1')
// (8, 3, 'lutff_0/in_2')
// (8, 3, 'lutff_2/in_3')
// (8, 3, 'lutff_4/in_1')
// (8, 3, 'lutff_5/in_2')
// (8, 3, 'sp4_r_v_b_33')
// (8, 4, 'neigh_op_top_4')
// (8, 4, 'sp4_r_v_b_20')
// (8, 5, 'lutff_4/out')
// (8, 5, 'sp4_r_v_b_9')
// (8, 6, 'neigh_op_bot_4')
// (9, 1, 'sp4_v_t_44')
// (9, 2, 'sp4_v_b_44')
// (9, 3, 'sp4_v_b_33')
// (9, 4, 'neigh_op_tnl_4')
// (9, 4, 'sp4_v_b_20')
// (9, 5, 'neigh_op_lft_4')
// (9, 5, 'sp4_v_b_9')
// (9, 6, 'neigh_op_bnl_4')

wire n431;
// (7, 4, 'neigh_op_tnr_5')
// (7, 5, 'neigh_op_rgt_5')
// (7, 6, 'neigh_op_bnr_5')
// (8, 4, 'local_g0_5')
// (8, 4, 'local_g1_5')
// (8, 4, 'lutff_3/in_0')
// (8, 4, 'lutff_6/in_1')
// (8, 4, 'lutff_7/in_1')
// (8, 4, 'neigh_op_top_5')
// (8, 5, 'lutff_5/out')
// (8, 6, 'neigh_op_bot_5')
// (9, 4, 'neigh_op_tnl_5')
// (9, 5, 'neigh_op_lft_5')
// (9, 6, 'neigh_op_bnl_5')

wire n432;
// (7, 4, 'neigh_op_tnr_6')
// (7, 5, 'neigh_op_rgt_6')
// (7, 6, 'neigh_op_bnr_6')
// (8, 0, 'span12_vert_20')
// (8, 1, 'sp12_v_b_20')
// (8, 2, 'sp12_v_b_19')
// (8, 3, 'local_g2_0')
// (8, 3, 'local_g3_0')
// (8, 3, 'lutff_0/in_1')
// (8, 3, 'lutff_2/in_2')
// (8, 3, 'lutff_5/in_1')
// (8, 3, 'lutff_7/in_2')
// (8, 3, 'sp12_v_b_16')
// (8, 4, 'neigh_op_top_6')
// (8, 4, 'sp12_v_b_15')
// (8, 5, 'lutff_6/out')
// (8, 5, 'sp12_v_b_12')
// (8, 6, 'neigh_op_bot_6')
// (8, 6, 'sp12_v_b_11')
// (8, 7, 'sp12_v_b_8')
// (8, 8, 'sp12_v_b_7')
// (8, 9, 'sp12_v_b_4')
// (8, 10, 'sp12_v_b_3')
// (8, 11, 'sp12_v_b_0')
// (9, 4, 'neigh_op_tnl_6')
// (9, 5, 'neigh_op_lft_6')
// (9, 6, 'neigh_op_bnl_6')

reg n433 = 0;
// (7, 4, 'neigh_op_tnr_7')
// (7, 5, 'neigh_op_rgt_7')
// (7, 6, 'neigh_op_bnr_7')
// (8, 4, 'neigh_op_top_7')
// (8, 5, 'local_g3_7')
// (8, 5, 'lutff_3/in_3')
// (8, 5, 'lutff_7/out')
// (8, 6, 'neigh_op_bot_7')
// (9, 4, 'neigh_op_tnl_7')
// (9, 5, 'neigh_op_lft_7')
// (9, 6, 'neigh_op_bnl_7')

wire n434;
// (7, 4, 'sp4_h_r_8')
// (8, 4, 'sp4_h_r_21')
// (9, 4, 'local_g2_0')
// (9, 4, 'local_g3_0')
// (9, 4, 'lutff_0/in_2')
// (9, 4, 'lutff_5/in_0')
// (9, 4, 'sp4_h_r_32')
// (10, 1, 'sp4_r_v_b_45')
// (10, 2, 'sp4_r_v_b_32')
// (10, 3, 'neigh_op_tnr_4')
// (10, 3, 'sp4_r_v_b_21')
// (10, 4, 'neigh_op_rgt_4')
// (10, 4, 'sp4_h_r_45')
// (10, 4, 'sp4_r_v_b_8')
// (10, 5, 'neigh_op_bnr_4')
// (11, 0, 'span4_vert_45')
// (11, 1, 'sp4_v_b_45')
// (11, 2, 'sp4_v_b_32')
// (11, 3, 'neigh_op_top_4')
// (11, 3, 'sp4_v_b_21')
// (11, 4, 'local_g3_4')
// (11, 4, 'lutff_4/out')
// (11, 4, 'lutff_7/in_0')
// (11, 4, 'sp4_h_l_45')
// (11, 4, 'sp4_v_b_8')
// (11, 5, 'neigh_op_bot_4')
// (12, 3, 'neigh_op_tnl_4')
// (12, 4, 'neigh_op_lft_4')
// (12, 5, 'neigh_op_bnl_4')

wire n435;
// (7, 4, 'sp4_r_v_b_46')
// (7, 5, 'neigh_op_tnr_3')
// (7, 5, 'sp4_r_v_b_35')
// (7, 6, 'neigh_op_rgt_3')
// (7, 6, 'sp4_r_v_b_22')
// (7, 7, 'neigh_op_bnr_3')
// (7, 7, 'sp4_r_v_b_11')
// (8, 3, 'sp4_v_t_46')
// (8, 4, 'sp4_v_b_46')
// (8, 5, 'local_g2_3')
// (8, 5, 'lutff_2/in_3')
// (8, 5, 'lutff_4/in_3')
// (8, 5, 'neigh_op_top_3')
// (8, 5, 'sp4_v_b_35')
// (8, 6, 'lutff_3/out')
// (8, 6, 'sp4_v_b_22')
// (8, 7, 'neigh_op_bot_3')
// (8, 7, 'sp4_v_b_11')
// (9, 5, 'neigh_op_tnl_3')
// (9, 6, 'neigh_op_lft_3')
// (9, 7, 'neigh_op_bnl_3')

wire n436;
// (7, 5, 'neigh_op_tnr_0')
// (7, 6, 'neigh_op_rgt_0')
// (7, 7, 'neigh_op_bnr_0')
// (8, 5, 'local_g0_0')
// (8, 5, 'lutff_2/in_2')
// (8, 5, 'neigh_op_top_0')
// (8, 6, 'lutff_0/out')
// (8, 7, 'neigh_op_bot_0')
// (9, 5, 'neigh_op_tnl_0')
// (9, 6, 'neigh_op_lft_0')
// (9, 7, 'neigh_op_bnl_0')

wire n437;
// (7, 5, 'neigh_op_tnr_1')
// (7, 6, 'neigh_op_rgt_1')
// (7, 7, 'neigh_op_bnr_1')
// (8, 3, 'sp4_r_v_b_38')
// (8, 4, 'local_g0_3')
// (8, 4, 'local_g1_3')
// (8, 4, 'lutff_0/in_2')
// (8, 4, 'lutff_1/in_2')
// (8, 4, 'sp4_r_v_b_27')
// (8, 5, 'neigh_op_top_1')
// (8, 5, 'sp4_r_v_b_14')
// (8, 6, 'lutff_1/out')
// (8, 6, 'sp4_r_v_b_3')
// (8, 7, 'neigh_op_bot_1')
// (9, 2, 'sp4_v_t_38')
// (9, 3, 'sp4_v_b_38')
// (9, 4, 'sp4_v_b_27')
// (9, 5, 'neigh_op_tnl_1')
// (9, 5, 'sp4_v_b_14')
// (9, 6, 'neigh_op_lft_1')
// (9, 6, 'sp4_v_b_3')
// (9, 7, 'neigh_op_bnl_1')

wire n438;
// (7, 5, 'neigh_op_tnr_2')
// (7, 6, 'neigh_op_rgt_2')
// (7, 7, 'neigh_op_bnr_2')
// (8, 0, 'span12_vert_15')
// (8, 1, 'sp12_v_b_15')
// (8, 2, 'sp12_v_b_12')
// (8, 3, 'sp12_v_b_11')
// (8, 4, 'local_g3_0')
// (8, 4, 'lutff_1/in_0')
// (8, 4, 'lutff_5/in_2')
// (8, 4, 'sp12_v_b_8')
// (8, 5, 'neigh_op_top_2')
// (8, 5, 'sp12_v_b_7')
// (8, 6, 'lutff_2/out')
// (8, 6, 'sp12_v_b_4')
// (8, 7, 'neigh_op_bot_2')
// (8, 7, 'sp12_v_b_3')
// (8, 8, 'sp12_v_b_0')
// (9, 5, 'neigh_op_tnl_2')
// (9, 6, 'neigh_op_lft_2')
// (9, 7, 'neigh_op_bnl_2')

wire n439;
// (7, 5, 'neigh_op_tnr_4')
// (7, 6, 'neigh_op_rgt_4')
// (7, 7, 'neigh_op_bnr_4')
// (8, 3, 'sp4_r_v_b_44')
// (8, 4, 'local_g0_2')
// (8, 4, 'local_g2_1')
// (8, 4, 'lutff_0/in_1')
// (8, 4, 'lutff_1/in_1')
// (8, 4, 'sp4_r_v_b_33')
// (8, 5, 'neigh_op_top_4')
// (8, 5, 'sp4_r_v_b_20')
// (8, 6, 'lutff_4/out')
// (8, 6, 'sp4_r_v_b_9')
// (8, 7, 'neigh_op_bot_4')
// (9, 2, 'sp4_v_t_44')
// (9, 3, 'sp4_v_b_44')
// (9, 4, 'sp4_v_b_33')
// (9, 5, 'neigh_op_tnl_4')
// (9, 5, 'sp4_v_b_20')
// (9, 6, 'neigh_op_lft_4')
// (9, 6, 'sp4_v_b_9')
// (9, 7, 'neigh_op_bnl_4')

reg n440 = 0;
// (7, 5, 'neigh_op_tnr_5')
// (7, 6, 'neigh_op_rgt_5')
// (7, 7, 'neigh_op_bnr_5')
// (8, 5, 'neigh_op_top_5')
// (8, 6, 'local_g1_5')
// (8, 6, 'lutff_3/in_3')
// (8, 6, 'lutff_5/out')
// (8, 7, 'neigh_op_bot_5')
// (9, 5, 'neigh_op_tnl_5')
// (9, 6, 'neigh_op_lft_5')
// (9, 7, 'neigh_op_bnl_5')

reg n441 = 0;
// (7, 5, 'neigh_op_tnr_6')
// (7, 6, 'neigh_op_rgt_6')
// (7, 7, 'neigh_op_bnr_6')
// (8, 5, 'neigh_op_top_6')
// (8, 6, 'local_g0_6')
// (8, 6, 'lutff_1/in_3')
// (8, 6, 'lutff_6/out')
// (8, 7, 'neigh_op_bot_6')
// (9, 5, 'neigh_op_tnl_6')
// (9, 6, 'neigh_op_lft_6')
// (9, 7, 'neigh_op_bnl_6')

reg n442 = 0;
// (7, 5, 'neigh_op_tnr_7')
// (7, 6, 'neigh_op_rgt_7')
// (7, 7, 'neigh_op_bnr_7')
// (8, 5, 'local_g0_7')
// (8, 5, 'lutff_0/in_3')
// (8, 5, 'neigh_op_top_7')
// (8, 6, 'lutff_7/out')
// (8, 7, 'neigh_op_bot_7')
// (9, 5, 'neigh_op_tnl_7')
// (9, 6, 'neigh_op_lft_7')
// (9, 7, 'neigh_op_bnl_7')

wire n443;
// (7, 6, 'neigh_op_tnr_0')
// (7, 7, 'neigh_op_rgt_0')
// (7, 8, 'neigh_op_bnr_0')
// (8, 6, 'neigh_op_top_0')
// (8, 7, 'local_g2_0')
// (8, 7, 'lutff_0/out')
// (8, 7, 'lutff_5/in_3')
// (8, 8, 'neigh_op_bot_0')
// (9, 6, 'neigh_op_tnl_0')
// (9, 7, 'neigh_op_lft_0')
// (9, 8, 'neigh_op_bnl_0')

wire n444;
// (7, 6, 'neigh_op_tnr_1')
// (7, 7, 'neigh_op_rgt_1')
// (7, 8, 'neigh_op_bnr_1')
// (8, 4, 'sp4_r_v_b_38')
// (8, 5, 'local_g0_3')
// (8, 5, 'local_g1_3')
// (8, 5, 'lutff_5/in_3')
// (8, 5, 'lutff_6/in_3')
// (8, 5, 'sp4_r_v_b_27')
// (8, 6, 'neigh_op_top_1')
// (8, 6, 'sp4_r_v_b_14')
// (8, 7, 'lutff_1/out')
// (8, 7, 'sp4_r_v_b_3')
// (8, 8, 'neigh_op_bot_1')
// (9, 3, 'sp4_v_t_38')
// (9, 4, 'sp4_v_b_38')
// (9, 5, 'sp4_v_b_27')
// (9, 6, 'neigh_op_tnl_1')
// (9, 6, 'sp4_v_b_14')
// (9, 7, 'neigh_op_lft_1')
// (9, 7, 'sp4_v_b_3')
// (9, 8, 'neigh_op_bnl_1')

wire n445;
// (7, 6, 'neigh_op_tnr_3')
// (7, 7, 'neigh_op_rgt_3')
// (7, 8, 'neigh_op_bnr_3')
// (8, 0, 'span12_vert_18')
// (8, 1, 'sp12_v_b_18')
// (8, 2, 'sp12_v_b_17')
// (8, 3, 'sp12_v_b_14')
// (8, 4, 'sp12_v_b_13')
// (8, 5, 'local_g3_2')
// (8, 5, 'lutff_2/in_1')
// (8, 5, 'sp12_v_b_10')
// (8, 6, 'neigh_op_top_3')
// (8, 6, 'sp12_v_b_9')
// (8, 7, 'lutff_3/out')
// (8, 7, 'sp12_v_b_6')
// (8, 8, 'neigh_op_bot_3')
// (8, 8, 'sp12_v_b_5')
// (8, 9, 'sp12_v_b_2')
// (8, 10, 'sp12_v_b_1')
// (9, 6, 'neigh_op_tnl_3')
// (9, 7, 'neigh_op_lft_3')
// (9, 8, 'neigh_op_bnl_3')

wire n446;
// (7, 6, 'neigh_op_tnr_4')
// (7, 7, 'neigh_op_rgt_4')
// (7, 8, 'neigh_op_bnr_4')
// (8, 4, 'sp4_r_v_b_44')
// (8, 5, 'local_g0_2')
// (8, 5, 'local_g2_1')
// (8, 5, 'lutff_5/in_2')
// (8, 5, 'lutff_6/in_0')
// (8, 5, 'sp4_r_v_b_33')
// (8, 6, 'neigh_op_top_4')
// (8, 6, 'sp4_r_v_b_20')
// (8, 7, 'lutff_4/out')
// (8, 7, 'sp4_r_v_b_9')
// (8, 8, 'neigh_op_bot_4')
// (9, 3, 'sp4_v_t_44')
// (9, 4, 'sp4_v_b_44')
// (9, 5, 'sp4_v_b_33')
// (9, 6, 'neigh_op_tnl_4')
// (9, 6, 'sp4_v_b_20')
// (9, 7, 'neigh_op_lft_4')
// (9, 7, 'sp4_v_b_9')
// (9, 8, 'neigh_op_bnl_4')

wire n447;
// (7, 6, 'neigh_op_tnr_5')
// (7, 7, 'neigh_op_rgt_5')
// (7, 8, 'neigh_op_bnr_5')
// (8, 0, 'span12_vert_22')
// (8, 1, 'sp12_v_b_22')
// (8, 2, 'sp12_v_b_21')
// (8, 3, 'local_g2_2')
// (8, 3, 'local_g3_2')
// (8, 3, 'lutff_0/in_3')
// (8, 3, 'lutff_4/in_2')
// (8, 3, 'sp12_v_b_18')
// (8, 4, 'sp12_v_b_17')
// (8, 5, 'sp12_v_b_14')
// (8, 6, 'neigh_op_top_5')
// (8, 6, 'sp12_v_b_13')
// (8, 7, 'lutff_5/out')
// (8, 7, 'sp12_v_b_10')
// (8, 8, 'neigh_op_bot_5')
// (8, 8, 'sp12_v_b_9')
// (8, 9, 'sp12_v_b_6')
// (8, 10, 'sp12_v_b_5')
// (8, 11, 'sp12_v_b_2')
// (8, 12, 'sp12_v_b_1')
// (9, 6, 'neigh_op_tnl_5')
// (9, 7, 'neigh_op_lft_5')
// (9, 8, 'neigh_op_bnl_5')

reg n448 = 0;
// (7, 6, 'neigh_op_tnr_6')
// (7, 7, 'neigh_op_rgt_6')
// (7, 8, 'neigh_op_bnr_6')
// (8, 6, 'neigh_op_top_6')
// (8, 7, 'local_g0_6')
// (8, 7, 'lutff_1/in_3')
// (8, 7, 'lutff_6/out')
// (8, 8, 'neigh_op_bot_6')
// (9, 6, 'neigh_op_tnl_6')
// (9, 7, 'neigh_op_lft_6')
// (9, 8, 'neigh_op_bnl_6')

reg n449 = 0;
// (7, 6, 'neigh_op_tnr_7')
// (7, 7, 'neigh_op_rgt_7')
// (7, 8, 'neigh_op_bnr_7')
// (8, 6, 'local_g0_7')
// (8, 6, 'lutff_0/in_3')
// (8, 6, 'neigh_op_top_7')
// (8, 7, 'lutff_7/out')
// (8, 8, 'neigh_op_bot_7')
// (9, 6, 'neigh_op_tnl_7')
// (9, 7, 'neigh_op_lft_7')
// (9, 8, 'neigh_op_bnl_7')

reg n450 = 0;
// (7, 7, 'neigh_op_tnr_3')
// (7, 8, 'neigh_op_rgt_3')
// (7, 9, 'neigh_op_bnr_3')
// (8, 7, 'local_g1_3')
// (8, 7, 'lutff_5/in_1')
// (8, 7, 'neigh_op_top_3')
// (8, 8, 'lutff_3/out')
// (8, 9, 'neigh_op_bot_3')
// (9, 7, 'neigh_op_tnl_3')
// (9, 8, 'neigh_op_lft_3')
// (9, 9, 'neigh_op_bnl_3')

reg n451 = 0;
// (7, 7, 'sp4_r_v_b_41')
// (7, 8, 'sp4_r_v_b_28')
// (7, 9, 'neigh_op_tnr_2')
// (7, 9, 'sp4_r_v_b_17')
// (7, 10, 'neigh_op_rgt_2')
// (7, 10, 'sp4_r_v_b_4')
// (7, 11, 'neigh_op_bnr_2')
// (8, 6, 'sp4_v_t_41')
// (8, 7, 'sp4_v_b_41')
// (8, 8, 'sp4_v_b_28')
// (8, 9, 'local_g1_1')
// (8, 9, 'lutff_2/in_0')
// (8, 9, 'neigh_op_top_2')
// (8, 9, 'sp4_v_b_17')
// (8, 10, 'local_g0_2')
// (8, 10, 'lutff_1/in_1')
// (8, 10, 'lutff_2/out')
// (8, 10, 'sp4_v_b_4')
// (8, 11, 'neigh_op_bot_2')
// (9, 9, 'neigh_op_tnl_2')
// (9, 10, 'neigh_op_lft_2')
// (9, 11, 'neigh_op_bnl_2')

wire n452;
// (7, 8, 'neigh_op_tnr_2')
// (7, 9, 'neigh_op_rgt_2')
// (7, 10, 'neigh_op_bnr_2')
// (8, 8, 'neigh_op_top_2')
// (8, 9, 'local_g2_2')
// (8, 9, 'lutff_1/in_3')
// (8, 9, 'lutff_2/out')
// (8, 10, 'neigh_op_bot_2')
// (9, 8, 'neigh_op_tnl_2')
// (9, 9, 'neigh_op_lft_2')
// (9, 10, 'neigh_op_bnl_2')

reg n453 = 0;
// (7, 8, 'neigh_op_tnr_3')
// (7, 9, 'neigh_op_rgt_3')
// (7, 10, 'neigh_op_bnr_3')
// (8, 8, 'neigh_op_top_3')
// (8, 9, 'local_g3_3')
// (8, 9, 'lutff_3/out')
// (8, 9, 'lutff_6/in_0')
// (8, 10, 'neigh_op_bot_3')
// (9, 8, 'neigh_op_tnl_3')
// (9, 9, 'neigh_op_lft_3')
// (9, 10, 'neigh_op_bnl_3')

reg n454 = 0;
// (7, 8, 'neigh_op_tnr_4')
// (7, 9, 'neigh_op_rgt_4')
// (7, 10, 'neigh_op_bnr_4')
// (8, 8, 'neigh_op_top_4')
// (8, 9, 'local_g0_4')
// (8, 9, 'local_g1_4')
// (8, 9, 'lutff_2/in_1')
// (8, 9, 'lutff_4/out')
// (8, 9, 'lutff_7/in_1')
// (8, 10, 'neigh_op_bot_4')
// (9, 8, 'neigh_op_tnl_4')
// (9, 9, 'neigh_op_lft_4')
// (9, 10, 'neigh_op_bnl_4')

reg n455 = 0;
// (7, 8, 'neigh_op_tnr_5')
// (7, 9, 'neigh_op_rgt_5')
// (7, 10, 'neigh_op_bnr_5')
// (8, 8, 'neigh_op_top_5')
// (8, 9, 'local_g1_5')
// (8, 9, 'lutff_4/in_0')
// (8, 9, 'lutff_5/out')
// (8, 10, 'neigh_op_bot_5')
// (9, 8, 'neigh_op_tnl_5')
// (9, 9, 'neigh_op_lft_5')
// (9, 10, 'neigh_op_bnl_5')

reg n456 = 0;
// (7, 8, 'neigh_op_tnr_6')
// (7, 9, 'neigh_op_rgt_6')
// (7, 10, 'neigh_op_bnr_6')
// (8, 8, 'neigh_op_top_6')
// (8, 9, 'local_g1_6')
// (8, 9, 'lutff_5/in_0')
// (8, 9, 'lutff_6/out')
// (8, 10, 'neigh_op_bot_6')
// (9, 8, 'neigh_op_tnl_6')
// (9, 9, 'neigh_op_lft_6')
// (9, 10, 'neigh_op_bnl_6')

reg n457 = 0;
// (7, 8, 'neigh_op_tnr_7')
// (7, 9, 'neigh_op_rgt_7')
// (7, 10, 'neigh_op_bnr_7')
// (8, 8, 'neigh_op_top_7')
// (8, 9, 'lutff_7/out')
// (8, 10, 'local_g1_7')
// (8, 10, 'lutff_0/in_0')
// (8, 10, 'neigh_op_bot_7')
// (9, 8, 'neigh_op_tnl_7')
// (9, 9, 'neigh_op_lft_7')
// (9, 10, 'neigh_op_bnl_7')

reg n458 = 0;
// (7, 9, 'neigh_op_tnr_0')
// (7, 10, 'neigh_op_rgt_0')
// (7, 11, 'neigh_op_bnr_0')
// (8, 9, 'neigh_op_top_0')
// (8, 10, 'local_g0_0')
// (8, 10, 'lutff_0/out')
// (8, 10, 'lutff_6/in_0')
// (8, 11, 'neigh_op_bot_0')
// (9, 9, 'neigh_op_tnl_0')
// (9, 10, 'neigh_op_lft_0')
// (9, 11, 'neigh_op_bnl_0')

reg n459 = 0;
// (7, 9, 'neigh_op_tnr_1')
// (7, 10, 'neigh_op_rgt_1')
// (7, 11, 'neigh_op_bnr_1')
// (8, 9, 'neigh_op_top_1')
// (8, 10, 'local_g0_1')
// (8, 10, 'lutff_1/out')
// (8, 10, 'lutff_7/in_0')
// (8, 11, 'neigh_op_bot_1')
// (9, 9, 'neigh_op_tnl_1')
// (9, 10, 'neigh_op_lft_1')
// (9, 11, 'neigh_op_bnl_1')

reg n460 = 0;
// (7, 9, 'neigh_op_tnr_3')
// (7, 10, 'neigh_op_rgt_3')
// (7, 11, 'neigh_op_bnr_3')
// (8, 9, 'neigh_op_top_3')
// (8, 10, 'local_g0_3')
// (8, 10, 'lutff_3/out')
// (8, 10, 'lutff_5/in_0')
// (8, 11, 'neigh_op_bot_3')
// (9, 9, 'neigh_op_tnl_3')
// (9, 10, 'neigh_op_lft_3')
// (9, 11, 'neigh_op_bnl_3')

reg n461 = 0;
// (7, 9, 'neigh_op_tnr_5')
// (7, 10, 'neigh_op_rgt_5')
// (7, 11, 'neigh_op_bnr_5')
// (8, 9, 'local_g0_5')
// (8, 9, 'lutff_1/in_0')
// (8, 9, 'lutff_3/in_0')
// (8, 9, 'lutff_7/in_0')
// (8, 9, 'neigh_op_top_5')
// (8, 10, 'local_g2_5')
// (8, 10, 'lutff_1/in_0')
// (8, 10, 'lutff_5/out')
// (8, 11, 'neigh_op_bot_5')
// (9, 9, 'neigh_op_tnl_5')
// (9, 10, 'neigh_op_lft_5')
// (9, 11, 'neigh_op_bnl_5')

reg n462 = 0;
// (7, 9, 'neigh_op_tnr_6')
// (7, 10, 'neigh_op_rgt_6')
// (7, 11, 'neigh_op_bnr_6')
// (8, 9, 'neigh_op_top_6')
// (8, 10, 'local_g0_6')
// (8, 10, 'lutff_2/in_0')
// (8, 10, 'lutff_6/out')
// (8, 11, 'neigh_op_bot_6')
// (9, 9, 'neigh_op_tnl_6')
// (9, 10, 'neigh_op_lft_6')
// (9, 11, 'neigh_op_bnl_6')

reg n463 = 0;
// (7, 9, 'neigh_op_tnr_7')
// (7, 10, 'neigh_op_rgt_7')
// (7, 11, 'neigh_op_bnr_7')
// (8, 9, 'neigh_op_top_7')
// (8, 10, 'local_g0_7')
// (8, 10, 'lutff_3/in_0')
// (8, 10, 'lutff_7/out')
// (8, 11, 'neigh_op_bot_7')
// (9, 9, 'neigh_op_tnl_7')
// (9, 10, 'neigh_op_lft_7')
// (9, 11, 'neigh_op_bnl_7')

reg n464 = 0;
// (7, 10, 'neigh_op_tnr_0')
// (7, 11, 'neigh_op_rgt_0')
// (7, 12, 'neigh_op_bnr_0')
// (8, 8, 'sp4_r_v_b_36')
// (8, 9, 'sp4_r_v_b_25')
// (8, 10, 'neigh_op_top_0')
// (8, 10, 'sp4_r_v_b_12')
// (8, 11, 'lutff_0/out')
// (8, 11, 'sp4_r_v_b_1')
// (8, 12, 'neigh_op_bot_0')
// (9, 7, 'sp4_v_t_36')
// (9, 8, 'sp4_v_b_36')
// (9, 9, 'sp4_v_b_25')
// (9, 10, 'neigh_op_tnl_0')
// (9, 10, 'sp4_v_b_12')
// (9, 11, 'local_g0_1')
// (9, 11, 'lutff_3/in_0')
// (9, 11, 'neigh_op_lft_0')
// (9, 11, 'sp4_v_b_1')
// (9, 12, 'neigh_op_bnl_0')

reg n465 = 0;
// (7, 10, 'neigh_op_tnr_1')
// (7, 11, 'neigh_op_rgt_1')
// (7, 12, 'neigh_op_bnr_1')
// (8, 10, 'neigh_op_top_1')
// (8, 11, 'local_g2_1')
// (8, 11, 'lutff_1/out')
// (8, 11, 'lutff_7/in_0')
// (8, 12, 'neigh_op_bot_1')
// (9, 10, 'neigh_op_tnl_1')
// (9, 11, 'neigh_op_lft_1')
// (9, 12, 'neigh_op_bnl_1')

reg n466 = 0;
// (7, 10, 'neigh_op_tnr_2')
// (7, 11, 'neigh_op_rgt_2')
// (7, 12, 'neigh_op_bnr_2')
// (8, 10, 'neigh_op_top_2')
// (8, 11, 'lutff_2/out')
// (8, 12, 'neigh_op_bot_2')
// (9, 10, 'neigh_op_tnl_2')
// (9, 11, 'local_g0_2')
// (9, 11, 'lutff_6/in_0')
// (9, 11, 'neigh_op_lft_2')
// (9, 12, 'neigh_op_bnl_2')

reg n467 = 0;
// (7, 10, 'neigh_op_tnr_3')
// (7, 11, 'neigh_op_rgt_3')
// (7, 12, 'neigh_op_bnr_3')
// (8, 10, 'neigh_op_top_3')
// (8, 11, 'local_g0_3')
// (8, 11, 'lutff_3/out')
// (8, 11, 'lutff_5/in_0')
// (8, 12, 'neigh_op_bot_3')
// (9, 10, 'neigh_op_tnl_3')
// (9, 11, 'neigh_op_lft_3')
// (9, 12, 'neigh_op_bnl_3')

reg n468 = 0;
// (7, 10, 'neigh_op_tnr_4')
// (7, 11, 'neigh_op_rgt_4')
// (7, 12, 'neigh_op_bnr_4')
// (8, 10, 'neigh_op_top_4')
// (8, 11, 'local_g1_4')
// (8, 11, 'lutff_1/in_0')
// (8, 11, 'lutff_4/out')
// (8, 12, 'neigh_op_bot_4')
// (9, 10, 'neigh_op_tnl_4')
// (9, 11, 'neigh_op_lft_4')
// (9, 12, 'neigh_op_bnl_4')

reg n469 = 0;
// (7, 10, 'neigh_op_tnr_5')
// (7, 11, 'neigh_op_rgt_5')
// (7, 12, 'neigh_op_bnr_5')
// (8, 10, 'neigh_op_top_5')
// (8, 11, 'lutff_5/out')
// (8, 12, 'local_g0_5')
// (8, 12, 'lutff_5/in_0')
// (8, 12, 'neigh_op_bot_5')
// (9, 10, 'neigh_op_tnl_5')
// (9, 11, 'neigh_op_lft_5')
// (9, 12, 'neigh_op_bnl_5')

reg n470 = 0;
// (7, 10, 'neigh_op_tnr_7')
// (7, 11, 'neigh_op_rgt_7')
// (7, 12, 'neigh_op_bnr_7')
// (8, 10, 'neigh_op_top_7')
// (8, 11, 'local_g1_7')
// (8, 11, 'lutff_0/in_0')
// (8, 11, 'lutff_7/out')
// (8, 12, 'neigh_op_bot_7')
// (9, 10, 'neigh_op_tnl_7')
// (9, 11, 'neigh_op_lft_7')
// (9, 12, 'neigh_op_bnl_7')

wire n471;
// (7, 11, 'local_g3_0')
// (7, 11, 'lutff_2/in_3')
// (7, 11, 'neigh_op_tnr_0')
// (7, 12, 'neigh_op_rgt_0')
// (7, 13, 'neigh_op_bnr_0')
// (8, 11, 'neigh_op_top_0')
// (8, 12, 'lutff_0/out')
// (8, 13, 'neigh_op_bot_0')
// (9, 11, 'neigh_op_tnl_0')
// (9, 12, 'neigh_op_lft_0')
// (9, 13, 'neigh_op_bnl_0')

reg n472 = 0;
// (7, 11, 'neigh_op_tnr_5')
// (7, 12, 'neigh_op_rgt_5')
// (7, 13, 'neigh_op_bnr_5')
// (8, 11, 'neigh_op_top_5')
// (8, 12, 'lutff_5/out')
// (8, 13, 'local_g1_5')
// (8, 13, 'lutff_4/in_0')
// (8, 13, 'neigh_op_bot_5')
// (9, 11, 'neigh_op_tnl_5')
// (9, 12, 'neigh_op_lft_5')
// (9, 13, 'neigh_op_bnl_5')

wire n473;
// (7, 12, 'neigh_op_tnr_1')
// (7, 13, 'neigh_op_rgt_1')
// (7, 14, 'neigh_op_bnr_1')
// (8, 11, 'sp4_r_v_b_43')
// (8, 12, 'local_g1_6')
// (8, 12, 'lutff_0/in_3')
// (8, 12, 'neigh_op_top_1')
// (8, 12, 'sp4_r_v_b_30')
// (8, 13, 'lutff_1/out')
// (8, 13, 'sp4_r_v_b_19')
// (8, 14, 'neigh_op_bot_1')
// (8, 14, 'sp4_r_v_b_6')
// (9, 10, 'sp4_v_t_43')
// (9, 11, 'sp4_v_b_43')
// (9, 12, 'neigh_op_tnl_1')
// (9, 12, 'sp4_v_b_30')
// (9, 13, 'neigh_op_lft_1')
// (9, 13, 'sp4_v_b_19')
// (9, 14, 'neigh_op_bnl_1')
// (9, 14, 'sp4_v_b_6')

reg n474 = 0;
// (7, 12, 'neigh_op_tnr_3')
// (7, 13, 'neigh_op_rgt_3')
// (7, 14, 'neigh_op_bnr_3')
// (8, 12, 'neigh_op_top_3')
// (8, 13, 'local_g0_3')
// (8, 13, 'local_g1_3')
// (8, 13, 'lutff_1/in_0')
// (8, 13, 'lutff_3/out')
// (8, 13, 'lutff_5/in_1')
// (8, 14, 'neigh_op_bot_3')
// (9, 12, 'neigh_op_tnl_3')
// (9, 13, 'neigh_op_lft_3')
// (9, 14, 'neigh_op_bnl_3')

reg n475 = 0;
// (7, 12, 'neigh_op_tnr_4')
// (7, 13, 'neigh_op_rgt_4')
// (7, 14, 'neigh_op_bnr_4')
// (8, 12, 'neigh_op_top_4')
// (8, 13, 'local_g0_4')
// (8, 13, 'local_g1_4')
// (8, 13, 'lutff_1/in_1')
// (8, 13, 'lutff_4/out')
// (8, 13, 'lutff_6/in_1')
// (8, 14, 'neigh_op_bot_4')
// (9, 12, 'neigh_op_tnl_4')
// (9, 13, 'neigh_op_lft_4')
// (9, 14, 'neigh_op_bnl_4')

reg n476 = 0;
// (7, 12, 'neigh_op_tnr_5')
// (7, 13, 'neigh_op_rgt_5')
// (7, 14, 'neigh_op_bnr_5')
// (8, 12, 'neigh_op_top_5')
// (8, 13, 'lutff_5/out')
// (8, 14, 'neigh_op_bot_5')
// (9, 12, 'neigh_op_tnl_5')
// (9, 13, 'local_g0_5')
// (9, 13, 'lutff_1/in_0')
// (9, 13, 'neigh_op_lft_5')
// (9, 14, 'neigh_op_bnl_5')

reg n477 = 0;
// (7, 12, 'neigh_op_tnr_6')
// (7, 13, 'neigh_op_rgt_6')
// (7, 14, 'neigh_op_bnr_6')
// (8, 12, 'neigh_op_top_6')
// (8, 13, 'local_g0_6')
// (8, 13, 'lutff_2/in_0')
// (8, 13, 'lutff_6/out')
// (8, 14, 'neigh_op_bot_6')
// (9, 12, 'neigh_op_tnl_6')
// (9, 13, 'neigh_op_lft_6')
// (9, 14, 'neigh_op_bnl_6')

reg n478 = 0;
// (7, 12, 'neigh_op_tnr_7')
// (7, 12, 'sp4_r_v_b_43')
// (7, 13, 'neigh_op_rgt_7')
// (7, 13, 'sp4_r_v_b_30')
// (7, 14, 'neigh_op_bnr_7')
// (7, 14, 'sp4_r_v_b_19')
// (7, 15, 'sp4_r_v_b_6')
// (8, 11, 'sp4_v_t_43')
// (8, 12, 'neigh_op_top_7')
// (8, 12, 'sp4_v_b_43')
// (8, 13, 'lutff_7/out')
// (8, 13, 'sp4_v_b_30')
// (8, 14, 'neigh_op_bot_7')
// (8, 14, 'sp4_v_b_19')
// (8, 15, 'local_g1_6')
// (8, 15, 'lutff_5/in_0')
// (8, 15, 'sp4_v_b_6')
// (9, 12, 'neigh_op_tnl_7')
// (9, 13, 'neigh_op_lft_7')
// (9, 14, 'neigh_op_bnl_7')

reg n479 = 0;
// (7, 13, 'neigh_op_tnr_0')
// (7, 14, 'neigh_op_rgt_0')
// (7, 15, 'neigh_op_bnr_0')
// (8, 13, 'neigh_op_top_0')
// (8, 14, 'local_g0_0')
// (8, 14, 'lutff_0/out')
// (8, 14, 'lutff_2/in_0')
// (8, 15, 'neigh_op_bot_0')
// (9, 13, 'neigh_op_tnl_0')
// (9, 14, 'neigh_op_lft_0')
// (9, 15, 'neigh_op_bnl_0')

reg n480 = 0;
// (7, 13, 'neigh_op_tnr_2')
// (7, 14, 'neigh_op_rgt_2')
// (7, 15, 'neigh_op_bnr_2')
// (8, 13, 'neigh_op_top_2')
// (8, 14, 'local_g0_2')
// (8, 14, 'lutff_2/out')
// (8, 14, 'lutff_6/in_0')
// (8, 15, 'neigh_op_bot_2')
// (9, 13, 'neigh_op_tnl_2')
// (9, 14, 'neigh_op_lft_2')
// (9, 15, 'neigh_op_bnl_2')

reg n481 = 0;
// (7, 13, 'neigh_op_tnr_6')
// (7, 14, 'neigh_op_rgt_6')
// (7, 15, 'neigh_op_bnr_6')
// (8, 8, 'sp12_v_t_23')
// (8, 9, 'sp12_v_b_23')
// (8, 10, 'sp12_v_b_20')
// (8, 11, 'local_g2_3')
// (8, 11, 'lutff_2/in_3')
// (8, 11, 'sp12_v_b_19')
// (8, 12, 'sp12_v_b_16')
// (8, 13, 'neigh_op_top_6')
// (8, 13, 'sp12_v_b_15')
// (8, 14, 'lutff_6/out')
// (8, 14, 'sp12_v_b_12')
// (8, 15, 'neigh_op_bot_6')
// (8, 15, 'sp12_v_b_11')
// (8, 16, 'sp12_v_b_8')
// (8, 17, 'span12_vert_7')
// (9, 13, 'neigh_op_tnl_6')
// (9, 14, 'neigh_op_lft_6')
// (9, 15, 'neigh_op_bnl_6')

reg n482 = 0;
// (7, 14, 'neigh_op_tnr_0')
// (7, 15, 'neigh_op_rgt_0')
// (7, 16, 'neigh_op_bnr_0')
// (8, 13, 'sp4_r_v_b_41')
// (8, 14, 'local_g0_4')
// (8, 14, 'lutff_0/in_0')
// (8, 14, 'neigh_op_top_0')
// (8, 14, 'sp4_r_v_b_28')
// (8, 15, 'lutff_0/out')
// (8, 15, 'sp4_r_v_b_17')
// (8, 16, 'neigh_op_bot_0')
// (8, 16, 'sp4_r_v_b_4')
// (9, 12, 'sp4_v_t_41')
// (9, 13, 'sp4_v_b_41')
// (9, 14, 'neigh_op_tnl_0')
// (9, 14, 'sp4_v_b_28')
// (9, 15, 'neigh_op_lft_0')
// (9, 15, 'sp4_v_b_17')
// (9, 16, 'neigh_op_bnl_0')
// (9, 16, 'sp4_v_b_4')

reg n483 = 0;
// (7, 14, 'neigh_op_tnr_2')
// (7, 15, 'neigh_op_rgt_2')
// (7, 16, 'neigh_op_bnr_2')
// (8, 14, 'neigh_op_top_2')
// (8, 15, 'local_g0_2')
// (8, 15, 'lutff_0/in_0')
// (8, 15, 'lutff_2/out')
// (8, 16, 'neigh_op_bot_2')
// (9, 14, 'neigh_op_tnl_2')
// (9, 15, 'neigh_op_lft_2')
// (9, 16, 'neigh_op_bnl_2')

reg n484 = 0;
// (7, 14, 'neigh_op_tnr_5')
// (7, 15, 'neigh_op_rgt_5')
// (7, 16, 'neigh_op_bnr_5')
// (8, 14, 'neigh_op_top_5')
// (8, 15, 'local_g1_5')
// (8, 15, 'lutff_5/out')
// (8, 15, 'lutff_6/in_0')
// (8, 16, 'neigh_op_bot_5')
// (9, 14, 'neigh_op_tnl_5')
// (9, 15, 'neigh_op_lft_5')
// (9, 16, 'neigh_op_bnl_5')

reg n485 = 0;
// (7, 14, 'neigh_op_tnr_6')
// (7, 15, 'neigh_op_rgt_6')
// (7, 16, 'neigh_op_bnr_6')
// (8, 14, 'neigh_op_top_6')
// (8, 15, 'local_g0_6')
// (8, 15, 'lutff_2/in_0')
// (8, 15, 'lutff_6/out')
// (8, 16, 'neigh_op_bot_6')
// (9, 14, 'neigh_op_tnl_6')
// (9, 15, 'neigh_op_lft_6')
// (9, 16, 'neigh_op_bnl_6')

wire n486;
// (8, 2, 'neigh_op_tnr_5')
// (8, 3, 'neigh_op_rgt_5')
// (8, 4, 'neigh_op_bnr_5')
// (9, 2, 'neigh_op_top_5')
// (9, 3, 'lutff_5/out')
// (9, 3, 'sp4_h_r_10')
// (9, 4, 'neigh_op_bot_5')
// (10, 2, 'neigh_op_tnl_5')
// (10, 3, 'neigh_op_lft_5')
// (10, 3, 'sp4_h_r_23')
// (10, 4, 'neigh_op_bnl_5')
// (11, 3, 'local_g2_2')
// (11, 3, 'lutff_global/cen')
// (11, 3, 'sp4_h_r_34')
// (12, 3, 'sp4_h_r_47')
// (13, 3, 'span4_horz_47')

wire n487;
// (8, 3, 'neigh_op_tnr_0')
// (8, 4, 'neigh_op_rgt_0')
// (8, 4, 'sp4_h_r_5')
// (8, 5, 'neigh_op_bnr_0')
// (9, 3, 'neigh_op_top_0')
// (9, 4, 'lutff_0/out')
// (9, 4, 'sp4_h_r_16')
// (9, 5, 'neigh_op_bot_0')
// (10, 3, 'neigh_op_tnl_0')
// (10, 4, 'neigh_op_lft_0')
// (10, 4, 'sp4_h_r_29')
// (10, 5, 'neigh_op_bnl_0')
// (11, 4, 'local_g2_0')
// (11, 4, 'lutff_1/in_3')
// (11, 4, 'sp4_h_r_40')
// (12, 4, 'sp4_h_l_40')

reg n488 = 0;
// (8, 3, 'neigh_op_tnr_4')
// (8, 4, 'neigh_op_rgt_4')
// (8, 5, 'neigh_op_bnr_4')
// (9, 3, 'neigh_op_top_4')
// (9, 4, 'local_g0_4')
// (9, 4, 'local_g1_4')
// (9, 4, 'lutff_0/in_1')
// (9, 4, 'lutff_4/in_1')
// (9, 4, 'lutff_4/out')
// (9, 4, 'lutff_7/in_3')
// (9, 4, 'sp4_h_r_8')
// (9, 4, 'sp4_r_v_b_41')
// (9, 5, 'neigh_op_bot_4')
// (9, 5, 'sp4_r_v_b_28')
// (9, 6, 'sp4_r_v_b_17')
// (9, 7, 'sp4_r_v_b_4')
// (10, 3, 'neigh_op_tnl_4')
// (10, 3, 'sp4_h_r_4')
// (10, 3, 'sp4_v_t_41')
// (10, 4, 'neigh_op_lft_4')
// (10, 4, 'sp4_h_r_21')
// (10, 4, 'sp4_v_b_41')
// (10, 5, 'neigh_op_bnl_4')
// (10, 5, 'sp4_v_b_28')
// (10, 6, 'sp4_v_b_17')
// (10, 7, 'sp4_v_b_4')
// (11, 3, 'local_g0_1')
// (11, 3, 'lutff_7/in_0')
// (11, 3, 'sp4_h_r_17')
// (11, 4, 'local_g3_0')
// (11, 4, 'lutff_6/in_3')
// (11, 4, 'sp4_h_r_32')
// (12, 3, 'sp4_h_r_28')
// (12, 4, 'sp4_h_r_45')
// (13, 3, 'span4_horz_28')
// (13, 4, 'span4_horz_45')

wire n489;
// (8, 4, 'neigh_op_tnr_1')
// (8, 5, 'neigh_op_rgt_1')
// (8, 6, 'neigh_op_bnr_1')
// (9, 4, 'neigh_op_top_1')
// (9, 5, 'lutff_1/out')
// (9, 6, 'local_g0_1')
// (9, 6, 'lutff_1/in_2')
// (9, 6, 'neigh_op_bot_1')
// (10, 4, 'neigh_op_tnl_1')
// (10, 5, 'neigh_op_lft_1')
// (10, 6, 'neigh_op_bnl_1')

reg n490 = 0;
// (8, 4, 'neigh_op_tnr_5')
// (8, 5, 'local_g3_5')
// (8, 5, 'lutff_1/in_3')
// (8, 5, 'neigh_op_rgt_5')
// (8, 6, 'neigh_op_bnr_5')
// (9, 4, 'neigh_op_top_5')
// (9, 5, 'lutff_5/out')
// (9, 6, 'local_g1_5')
// (9, 6, 'lutff_0/in_0')
// (9, 6, 'neigh_op_bot_5')
// (10, 4, 'neigh_op_tnl_5')
// (10, 5, 'neigh_op_lft_5')
// (10, 6, 'neigh_op_bnl_5')

reg n491 = 0;
// (8, 4, 'neigh_op_tnr_7')
// (8, 5, 'neigh_op_rgt_7')
// (8, 6, 'neigh_op_bnr_7')
// (9, 4, 'neigh_op_top_7')
// (9, 5, 'local_g0_7')
// (9, 5, 'lutff_5/in_0')
// (9, 5, 'lutff_7/out')
// (9, 6, 'neigh_op_bot_7')
// (10, 4, 'neigh_op_tnl_7')
// (10, 5, 'neigh_op_lft_7')
// (10, 6, 'neigh_op_bnl_7')

wire n492;
// (8, 4, 'sp4_h_r_7')
// (8, 5, 'sp4_h_r_3')
// (9, 4, 'local_g0_2')
// (9, 4, 'lutff_2/in_2')
// (9, 4, 'sp4_h_r_18')
// (9, 5, 'local_g1_6')
// (9, 5, 'lutff_1/in_2')
// (9, 5, 'sp4_h_r_14')
// (10, 3, 'neigh_op_tnr_3')
// (10, 4, 'neigh_op_rgt_3')
// (10, 4, 'sp4_h_r_31')
// (10, 5, 'neigh_op_bnr_3')
// (10, 5, 'sp4_h_r_27')
// (11, 1, 'sp4_r_v_b_42')
// (11, 2, 'sp4_r_v_b_31')
// (11, 2, 'sp4_r_v_b_47')
// (11, 3, 'neigh_op_top_3')
// (11, 3, 'sp4_r_v_b_18')
// (11, 3, 'sp4_r_v_b_34')
// (11, 4, 'lutff_3/out')
// (11, 4, 'sp4_h_r_42')
// (11, 4, 'sp4_r_v_b_23')
// (11, 4, 'sp4_r_v_b_7')
// (11, 5, 'neigh_op_bot_3')
// (11, 5, 'sp4_h_r_38')
// (11, 5, 'sp4_r_v_b_10')
// (12, 0, 'span4_vert_42')
// (12, 1, 'sp4_v_b_42')
// (12, 1, 'sp4_v_t_47')
// (12, 2, 'sp4_v_b_31')
// (12, 2, 'sp4_v_b_47')
// (12, 3, 'neigh_op_tnl_3')
// (12, 3, 'sp4_v_b_18')
// (12, 3, 'sp4_v_b_34')
// (12, 4, 'neigh_op_lft_3')
// (12, 4, 'sp4_h_l_42')
// (12, 4, 'sp4_v_b_23')
// (12, 4, 'sp4_v_b_7')
// (12, 5, 'neigh_op_bnl_3')
// (12, 5, 'sp4_h_l_38')
// (12, 5, 'sp4_v_b_10')

reg n493 = 0;
// (8, 4, 'sp4_r_v_b_41')
// (8, 5, 'sp4_r_v_b_28')
// (8, 6, 'neigh_op_tnr_2')
// (8, 6, 'sp4_r_v_b_17')
// (8, 7, 'neigh_op_rgt_2')
// (8, 7, 'sp4_r_v_b_4')
// (8, 8, 'neigh_op_bnr_2')
// (9, 3, 'sp4_v_t_41')
// (9, 4, 'local_g3_1')
// (9, 4, 'lutff_1/in_3')
// (9, 4, 'sp4_v_b_41')
// (9, 5, 'sp4_v_b_28')
// (9, 6, 'local_g0_2')
// (9, 6, 'lutff_6/in_0')
// (9, 6, 'neigh_op_top_2')
// (9, 6, 'sp4_v_b_17')
// (9, 7, 'lutff_2/out')
// (9, 7, 'sp4_v_b_4')
// (9, 8, 'neigh_op_bot_2')
// (10, 6, 'neigh_op_tnl_2')
// (10, 7, 'neigh_op_lft_2')
// (10, 8, 'neigh_op_bnl_2')

reg n494 = 0;
// (8, 5, 'neigh_op_tnr_4')
// (8, 6, 'neigh_op_rgt_4')
// (8, 7, 'neigh_op_bnr_4')
// (9, 5, 'neigh_op_top_4')
// (9, 6, 'local_g1_4')
// (9, 6, 'lutff_4/out')
// (9, 6, 'lutff_5/in_0')
// (9, 7, 'neigh_op_bot_4')
// (10, 5, 'neigh_op_tnl_4')
// (10, 6, 'neigh_op_lft_4')
// (10, 7, 'neigh_op_bnl_4')

reg n495 = 0;
// (8, 5, 'neigh_op_tnr_5')
// (8, 6, 'local_g2_5')
// (8, 6, 'lutff_2/in_3')
// (8, 6, 'neigh_op_rgt_5')
// (8, 7, 'neigh_op_bnr_5')
// (9, 5, 'neigh_op_top_5')
// (9, 6, 'local_g0_5')
// (9, 6, 'lutff_3/in_0')
// (9, 6, 'lutff_5/out')
// (9, 7, 'neigh_op_bot_5')
// (10, 5, 'neigh_op_tnl_5')
// (10, 6, 'neigh_op_lft_5')
// (10, 7, 'neigh_op_bnl_5')

reg n496 = 0;
// (8, 6, 'neigh_op_tnr_1')
// (8, 7, 'neigh_op_rgt_1')
// (8, 8, 'neigh_op_bnr_1')
// (9, 6, 'neigh_op_top_1')
// (9, 7, 'local_g0_1')
// (9, 7, 'lutff_1/out')
// (9, 7, 'lutff_7/in_0')
// (9, 8, 'neigh_op_bot_1')
// (10, 6, 'neigh_op_tnl_1')
// (10, 7, 'neigh_op_lft_1')
// (10, 8, 'neigh_op_bnl_1')

reg n497 = 0;
// (8, 6, 'neigh_op_tnr_3')
// (8, 7, 'neigh_op_rgt_3')
// (8, 8, 'neigh_op_bnr_3')
// (9, 6, 'neigh_op_top_3')
// (9, 7, 'local_g0_3')
// (9, 7, 'lutff_1/in_0')
// (9, 7, 'lutff_3/out')
// (9, 8, 'neigh_op_bot_3')
// (10, 6, 'neigh_op_tnl_3')
// (10, 7, 'neigh_op_lft_3')
// (10, 8, 'neigh_op_bnl_3')

reg n498 = 0;
// (8, 6, 'neigh_op_tnr_7')
// (8, 7, 'neigh_op_rgt_7')
// (8, 8, 'neigh_op_bnr_7')
// (9, 6, 'neigh_op_top_7')
// (9, 7, 'local_g1_7')
// (9, 7, 'lutff_0/in_0')
// (9, 7, 'lutff_7/out')
// (9, 8, 'neigh_op_bot_7')
// (10, 6, 'neigh_op_tnl_7')
// (10, 7, 'neigh_op_lft_7')
// (10, 8, 'neigh_op_bnl_7')

reg n499 = 0;
// (8, 7, 'neigh_op_tnr_3')
// (8, 8, 'neigh_op_rgt_3')
// (8, 8, 'sp4_h_r_11')
// (8, 9, 'neigh_op_bnr_3')
// (9, 7, 'neigh_op_top_3')
// (9, 8, 'lutff_3/out')
// (9, 8, 'sp4_h_r_22')
// (9, 9, 'neigh_op_bot_3')
// (10, 7, 'neigh_op_tnl_3')
// (10, 8, 'neigh_op_lft_3')
// (10, 8, 'sp4_h_r_35')
// (10, 9, 'neigh_op_bnl_3')
// (11, 8, 'sp4_h_r_46')
// (11, 9, 'sp4_r_v_b_41')
// (11, 10, 'local_g1_4')
// (11, 10, 'lutff_5/in_2')
// (11, 10, 'sp4_r_v_b_28')
// (11, 11, 'sp4_r_v_b_17')
// (11, 12, 'sp4_r_v_b_4')
// (12, 8, 'sp4_h_l_46')
// (12, 8, 'sp4_v_t_41')
// (12, 9, 'sp4_v_b_41')
// (12, 10, 'sp4_v_b_28')
// (12, 11, 'sp4_v_b_17')
// (12, 12, 'sp4_v_b_4')

reg n500 = 0;
// (8, 7, 'neigh_op_tnr_6')
// (8, 8, 'neigh_op_rgt_6')
// (8, 9, 'neigh_op_bnr_6')
// (9, 6, 'sp4_r_v_b_37')
// (9, 7, 'neigh_op_top_6')
// (9, 7, 'sp4_r_v_b_24')
// (9, 8, 'lutff_6/out')
// (9, 8, 'sp4_r_v_b_13')
// (9, 9, 'neigh_op_bot_6')
// (9, 9, 'sp4_r_v_b_0')
// (10, 5, 'sp4_v_t_37')
// (10, 6, 'sp4_v_b_37')
// (10, 7, 'neigh_op_tnl_6')
// (10, 7, 'sp4_v_b_24')
// (10, 8, 'neigh_op_lft_6')
// (10, 8, 'sp4_v_b_13')
// (10, 9, 'neigh_op_bnl_6')
// (10, 9, 'sp4_h_r_6')
// (10, 9, 'sp4_v_b_0')
// (11, 9, 'local_g0_3')
// (11, 9, 'lutff_3/in_0')
// (11, 9, 'sp4_h_r_19')
// (12, 9, 'sp4_h_r_30')
// (13, 9, 'span4_horz_30')

reg n501 = 0;
// (8, 8, 'neigh_op_tnr_0')
// (8, 9, 'neigh_op_rgt_0')
// (8, 10, 'neigh_op_bnr_0')
// (9, 8, 'neigh_op_top_0')
// (9, 9, 'local_g2_0')
// (9, 9, 'lutff_0/out')
// (9, 9, 'lutff_2/in_0')
// (9, 10, 'neigh_op_bot_0')
// (10, 8, 'neigh_op_tnl_0')
// (10, 9, 'neigh_op_lft_0')
// (10, 10, 'neigh_op_bnl_0')

reg n502 = 0;
// (8, 8, 'neigh_op_tnr_1')
// (8, 9, 'neigh_op_rgt_1')
// (8, 10, 'neigh_op_bnr_1')
// (9, 8, 'neigh_op_top_1')
// (9, 9, 'local_g1_1')
// (9, 9, 'lutff_0/in_0')
// (9, 9, 'lutff_1/out')
// (9, 10, 'neigh_op_bot_1')
// (10, 8, 'neigh_op_tnl_1')
// (10, 9, 'neigh_op_lft_1')
// (10, 10, 'neigh_op_bnl_1')

reg n503 = 0;
// (8, 8, 'neigh_op_tnr_2')
// (8, 9, 'neigh_op_rgt_2')
// (8, 9, 'sp4_h_r_9')
// (8, 10, 'neigh_op_bnr_2')
// (9, 8, 'neigh_op_top_2')
// (9, 9, 'lutff_2/out')
// (9, 9, 'sp4_h_r_20')
// (9, 10, 'neigh_op_bot_2')
// (10, 8, 'neigh_op_tnl_2')
// (10, 9, 'neigh_op_lft_2')
// (10, 9, 'sp4_h_r_33')
// (10, 10, 'neigh_op_bnl_2')
// (11, 9, 'local_g2_4')
// (11, 9, 'lutff_2/in_0')
// (11, 9, 'sp4_h_r_44')
// (12, 9, 'sp4_h_l_44')

reg n504 = 0;
// (8, 8, 'neigh_op_tnr_3')
// (8, 9, 'neigh_op_rgt_3')
// (8, 10, 'neigh_op_bnr_3')
// (9, 8, 'neigh_op_top_3')
// (9, 9, 'local_g1_3')
// (9, 9, 'lutff_3/out')
// (9, 9, 'lutff_7/in_3')
// (9, 10, 'neigh_op_bot_3')
// (10, 8, 'neigh_op_tnl_3')
// (10, 9, 'neigh_op_lft_3')
// (10, 10, 'neigh_op_bnl_3')

reg n505 = 0;
// (8, 8, 'neigh_op_tnr_4')
// (8, 9, 'neigh_op_rgt_4')
// (8, 10, 'neigh_op_bnr_4')
// (9, 8, 'neigh_op_top_4')
// (9, 9, 'local_g0_4')
// (9, 9, 'lutff_1/in_3')
// (9, 9, 'lutff_4/out')
// (9, 10, 'neigh_op_bot_4')
// (10, 8, 'neigh_op_tnl_4')
// (10, 9, 'neigh_op_lft_4')
// (10, 10, 'neigh_op_bnl_4')

reg n506 = 0;
// (8, 8, 'neigh_op_tnr_5')
// (8, 9, 'neigh_op_rgt_5')
// (8, 10, 'neigh_op_bnr_5')
// (9, 8, 'neigh_op_top_5')
// (9, 9, 'lutff_5/out')
// (9, 10, 'local_g1_5')
// (9, 10, 'lutff_0/in_0')
// (9, 10, 'neigh_op_bot_5')
// (10, 8, 'neigh_op_tnl_5')
// (10, 9, 'neigh_op_lft_5')
// (10, 10, 'neigh_op_bnl_5')

reg n507 = 0;
// (8, 8, 'neigh_op_tnr_6')
// (8, 9, 'neigh_op_rgt_6')
// (8, 10, 'neigh_op_bnr_6')
// (9, 8, 'neigh_op_top_6')
// (9, 9, 'local_g0_6')
// (9, 9, 'lutff_4/in_0')
// (9, 9, 'lutff_6/out')
// (9, 10, 'neigh_op_bot_6')
// (10, 8, 'neigh_op_tnl_6')
// (10, 9, 'neigh_op_lft_6')
// (10, 10, 'neigh_op_bnl_6')

reg n508 = 0;
// (8, 9, 'neigh_op_tnr_0')
// (8, 10, 'neigh_op_rgt_0')
// (8, 11, 'neigh_op_bnr_0')
// (9, 9, 'neigh_op_top_0')
// (9, 10, 'local_g1_0')
// (9, 10, 'lutff_0/out')
// (9, 10, 'lutff_7/in_0')
// (9, 11, 'neigh_op_bot_0')
// (10, 9, 'neigh_op_tnl_0')
// (10, 10, 'neigh_op_lft_0')
// (10, 11, 'neigh_op_bnl_0')

reg n509 = 0;
// (8, 9, 'neigh_op_tnr_2')
// (8, 10, 'neigh_op_rgt_2')
// (8, 11, 'neigh_op_bnr_2')
// (9, 9, 'local_g0_2')
// (9, 9, 'lutff_6/in_0')
// (9, 9, 'neigh_op_top_2')
// (9, 10, 'lutff_2/out')
// (9, 11, 'neigh_op_bot_2')
// (10, 9, 'neigh_op_tnl_2')
// (10, 10, 'neigh_op_lft_2')
// (10, 11, 'neigh_op_bnl_2')

reg n510 = 0;
// (8, 9, 'neigh_op_tnr_3')
// (8, 10, 'neigh_op_rgt_3')
// (8, 11, 'neigh_op_bnr_3')
// (9, 9, 'local_g0_3')
// (9, 9, 'lutff_3/in_0')
// (9, 9, 'neigh_op_top_3')
// (9, 10, 'lutff_3/out')
// (9, 11, 'neigh_op_bot_3')
// (10, 9, 'neigh_op_tnl_3')
// (10, 10, 'neigh_op_lft_3')
// (10, 11, 'neigh_op_bnl_3')

reg n511 = 0;
// (8, 9, 'neigh_op_tnr_5')
// (8, 10, 'neigh_op_rgt_5')
// (8, 11, 'neigh_op_bnr_5')
// (9, 9, 'neigh_op_top_5')
// (9, 10, 'local_g3_5')
// (9, 10, 'lutff_2/in_0')
// (9, 10, 'lutff_5/out')
// (9, 11, 'neigh_op_bot_5')
// (10, 9, 'neigh_op_tnl_5')
// (10, 10, 'neigh_op_lft_5')
// (10, 11, 'neigh_op_bnl_5')

reg n512 = 0;
// (8, 9, 'neigh_op_tnr_6')
// (8, 10, 'neigh_op_rgt_6')
// (8, 11, 'neigh_op_bnr_6')
// (9, 9, 'neigh_op_top_6')
// (9, 10, 'local_g1_6')
// (9, 10, 'lutff_5/in_0')
// (9, 10, 'lutff_6/out')
// (9, 11, 'neigh_op_bot_6')
// (10, 9, 'neigh_op_tnl_6')
// (10, 10, 'neigh_op_lft_6')
// (10, 11, 'neigh_op_bnl_6')

reg n513 = 0;
// (8, 9, 'neigh_op_tnr_7')
// (8, 10, 'neigh_op_rgt_7')
// (8, 11, 'neigh_op_bnr_7')
// (9, 9, 'neigh_op_top_7')
// (9, 10, 'local_g1_7')
// (9, 10, 'lutff_6/in_0')
// (9, 10, 'lutff_7/out')
// (9, 11, 'neigh_op_bot_7')
// (10, 9, 'neigh_op_tnl_7')
// (10, 10, 'neigh_op_lft_7')
// (10, 11, 'neigh_op_bnl_7')

wire \d_out[3] ;
// (8, 10, 'neigh_op_tnr_0')
// (8, 11, 'neigh_op_rgt_0')
// (8, 12, 'neigh_op_bnr_0')
// (9, 10, 'neigh_op_top_0')
// (9, 11, 'lutff_0/out')
// (9, 11, 'sp4_h_r_0')
// (9, 12, 'neigh_op_bot_0')
// (10, 10, 'neigh_op_tnl_0')
// (10, 11, 'neigh_op_lft_0')
// (10, 11, 'sp4_h_r_13')
// (10, 12, 'neigh_op_bnl_0')
// (11, 11, 'sp4_h_r_24')
// (12, 11, 'sp4_h_r_37')
// (13, 11, 'io_0/D_OUT_0')
// (13, 11, 'io_0/PAD')
// (13, 11, 'local_g1_5')
// (13, 11, 'span4_horz_37')

wire \d_out[0] ;
// (8, 10, 'neigh_op_tnr_1')
// (8, 11, 'neigh_op_rgt_1')
// (8, 12, 'neigh_op_bnr_1')
// (9, 9, 'sp4_r_v_b_43')
// (9, 10, 'neigh_op_top_1')
// (9, 10, 'sp4_r_v_b_30')
// (9, 11, 'lutff_1/out')
// (9, 11, 'sp4_r_v_b_19')
// (9, 12, 'neigh_op_bot_1')
// (9, 12, 'sp4_r_v_b_6')
// (10, 8, 'sp4_v_t_43')
// (10, 9, 'sp4_v_b_43')
// (10, 10, 'neigh_op_tnl_1')
// (10, 10, 'sp4_v_b_30')
// (10, 11, 'neigh_op_lft_1')
// (10, 11, 'sp4_v_b_19')
// (10, 12, 'neigh_op_bnl_1')
// (10, 12, 'sp4_h_r_0')
// (10, 12, 'sp4_v_b_6')
// (11, 12, 'sp4_h_r_13')
// (12, 12, 'sp4_h_r_24')
// (13, 12, 'io_1/D_OUT_0')
// (13, 12, 'io_1/PAD')
// (13, 12, 'local_g1_0')
// (13, 12, 'span4_horz_24')

reg n516 = 0;
// (8, 10, 'neigh_op_tnr_3')
// (8, 11, 'neigh_op_rgt_3')
// (8, 12, 'neigh_op_bnr_3')
// (9, 10, 'neigh_op_top_3')
// (9, 11, 'local_g1_3')
// (9, 11, 'lutff_3/out')
// (9, 11, 'lutff_4/in_0')
// (9, 12, 'neigh_op_bot_3')
// (10, 10, 'neigh_op_tnl_3')
// (10, 11, 'neigh_op_lft_3')
// (10, 12, 'neigh_op_bnl_3')

reg n517 = 0;
// (8, 10, 'neigh_op_tnr_4')
// (8, 11, 'neigh_op_rgt_4')
// (8, 12, 'neigh_op_bnr_4')
// (9, 10, 'local_g1_4')
// (9, 10, 'lutff_3/in_0')
// (9, 10, 'neigh_op_top_4')
// (9, 11, 'lutff_4/out')
// (9, 12, 'neigh_op_bot_4')
// (10, 10, 'neigh_op_tnl_4')
// (10, 11, 'neigh_op_lft_4')
// (10, 12, 'neigh_op_bnl_4')

reg n518 = 0;
// (8, 10, 'neigh_op_tnr_5')
// (8, 11, 'neigh_op_rgt_5')
// (8, 11, 'sp12_h_r_1')
// (8, 12, 'neigh_op_bnr_5')
// (9, 10, 'neigh_op_top_5')
// (9, 11, 'lutff_5/out')
// (9, 11, 'sp12_h_r_2')
// (9, 12, 'neigh_op_bot_5')
// (10, 10, 'neigh_op_tnl_5')
// (10, 11, 'neigh_op_lft_5')
// (10, 11, 'sp12_h_r_5')
// (10, 12, 'neigh_op_bnl_5')
// (11, 11, 'local_g1_6')
// (11, 11, 'lutff_3/in_0')
// (11, 11, 'sp12_h_r_6')
// (12, 11, 'sp12_h_r_9')
// (13, 11, 'span12_horz_9')

reg n519 = 0;
// (8, 10, 'neigh_op_tnr_6')
// (8, 11, 'neigh_op_rgt_6')
// (8, 12, 'neigh_op_bnr_6')
// (9, 10, 'neigh_op_top_6')
// (9, 11, 'local_g1_6')
// (9, 11, 'lutff_5/in_0')
// (9, 11, 'lutff_6/out')
// (9, 12, 'neigh_op_bot_6')
// (10, 10, 'neigh_op_tnl_6')
// (10, 11, 'neigh_op_lft_6')
// (10, 12, 'neigh_op_bnl_6')

wire \d_out[2] ;
// (8, 10, 'sp4_h_r_7')
// (9, 10, 'sp4_h_r_18')
// (10, 9, 'neigh_op_tnr_5')
// (10, 10, 'neigh_op_rgt_5')
// (10, 10, 'sp4_h_r_31')
// (10, 11, 'neigh_op_bnr_5')
// (11, 9, 'neigh_op_top_5')
// (11, 10, 'lutff_5/out')
// (11, 10, 'sp4_h_r_42')
// (11, 11, 'neigh_op_bot_5')
// (12, 9, 'neigh_op_tnl_5')
// (12, 10, 'neigh_op_lft_5')
// (12, 10, 'sp4_h_l_42')
// (12, 10, 'sp4_h_r_7')
// (12, 11, 'neigh_op_bnl_5')
// (13, 10, 'span4_horz_7')
// (13, 10, 'span4_vert_t_13')
// (13, 11, 'io_1/D_OUT_0')
// (13, 11, 'io_1/PAD')
// (13, 11, 'local_g0_5')
// (13, 11, 'span4_vert_b_13')
// (13, 12, 'span4_vert_b_9')
// (13, 13, 'span4_vert_b_5')
// (13, 14, 'span4_vert_b_1')

reg n521 = 0;
// (8, 10, 'sp4_r_v_b_36')
// (8, 11, 'local_g0_1')
// (8, 11, 'lutff_3/in_0')
// (8, 11, 'sp4_r_v_b_25')
// (8, 12, 'local_g2_4')
// (8, 12, 'lutff_0/in_0')
// (8, 12, 'neigh_op_tnr_4')
// (8, 12, 'sp4_r_v_b_12')
// (8, 13, 'local_g2_4')
// (8, 13, 'local_g3_4')
// (8, 13, 'lutff_5/in_0')
// (8, 13, 'lutff_6/in_0')
// (8, 13, 'neigh_op_rgt_4')
// (8, 13, 'sp4_r_v_b_1')
// (8, 14, 'neigh_op_bnr_4')
// (9, 9, 'sp4_v_t_36')
// (9, 10, 'sp4_v_b_36')
// (9, 11, 'sp4_v_b_25')
// (9, 12, 'neigh_op_top_4')
// (9, 12, 'sp4_v_b_12')
// (9, 13, 'lutff_4/out')
// (9, 13, 'sp4_h_r_8')
// (9, 13, 'sp4_v_b_1')
// (9, 14, 'neigh_op_bot_4')
// (10, 12, 'neigh_op_tnl_4')
// (10, 13, 'neigh_op_lft_4')
// (10, 13, 'sp4_h_r_21')
// (10, 14, 'neigh_op_bnl_4')
// (11, 13, 'sp4_h_r_32')
// (12, 13, 'sp4_h_r_45')
// (13, 13, 'span4_horz_45')

reg n522 = 0;
// (8, 11, 'neigh_op_tnr_4')
// (8, 12, 'neigh_op_rgt_4')
// (8, 13, 'neigh_op_bnr_4')
// (9, 11, 'neigh_op_top_4')
// (9, 12, 'local_g1_4')
// (9, 12, 'lutff_4/out')
// (9, 12, 'lutff_5/in_0')
// (9, 13, 'neigh_op_bot_4')
// (10, 11, 'neigh_op_tnl_4')
// (10, 12, 'neigh_op_lft_4')
// (10, 13, 'neigh_op_bnl_4')

reg n523 = 0;
// (8, 11, 'neigh_op_tnr_5')
// (8, 12, 'neigh_op_rgt_5')
// (8, 13, 'neigh_op_bnr_5')
// (9, 11, 'neigh_op_top_5')
// (9, 12, 'local_g1_5')
// (9, 12, 'lutff_2/in_0')
// (9, 12, 'lutff_5/out')
// (9, 13, 'neigh_op_bot_5')
// (10, 11, 'neigh_op_tnl_5')
// (10, 12, 'neigh_op_lft_5')
// (10, 13, 'neigh_op_bnl_5')

reg n524 = 0;
// (8, 12, 'neigh_op_tnr_1')
// (8, 13, 'neigh_op_rgt_1')
// (8, 14, 'neigh_op_bnr_1')
// (9, 12, 'neigh_op_top_1')
// (9, 13, 'local_g1_1')
// (9, 13, 'lutff_1/out')
// (9, 13, 'lutff_6/in_0')
// (9, 14, 'neigh_op_bot_1')
// (10, 12, 'neigh_op_tnl_1')
// (10, 13, 'neigh_op_lft_1')
// (10, 14, 'neigh_op_bnl_1')

reg n525 = 0;
// (8, 12, 'neigh_op_tnr_6')
// (8, 13, 'neigh_op_rgt_6')
// (8, 14, 'neigh_op_bnr_6')
// (9, 12, 'neigh_op_top_6')
// (9, 13, 'local_g0_6')
// (9, 13, 'lutff_4/in_0')
// (9, 13, 'lutff_6/out')
// (9, 14, 'neigh_op_bot_6')
// (10, 12, 'neigh_op_tnl_6')
// (10, 13, 'neigh_op_lft_6')
// (10, 14, 'neigh_op_bnl_6')

reg n526 = 0;
// (8, 13, 'local_g0_5')
// (8, 13, 'lutff_3/in_0')
// (8, 13, 'sp4_h_r_5')
// (9, 13, 'sp4_h_r_16')
// (10, 12, 'neigh_op_tnr_4')
// (10, 13, 'neigh_op_rgt_4')
// (10, 13, 'sp4_h_r_29')
// (10, 14, 'neigh_op_bnr_4')
// (11, 12, 'neigh_op_top_4')
// (11, 13, 'lutff_4/out')
// (11, 13, 'sp4_h_r_40')
// (11, 14, 'neigh_op_bot_4')
// (12, 12, 'neigh_op_tnl_4')
// (12, 13, 'neigh_op_lft_4')
// (12, 13, 'sp4_h_l_40')
// (12, 14, 'neigh_op_bnl_4')

wire n527;
// (9, 4, 'local_g0_0')
// (9, 4, 'local_g1_0')
// (9, 4, 'lutff_0/in_0')
// (9, 4, 'lutff_4/in_0')
// (9, 4, 'lutff_7/in_2')
// (9, 4, 'sp4_h_r_0')
// (10, 3, 'neigh_op_tnr_0')
// (10, 4, 'neigh_op_rgt_0')
// (10, 4, 'sp4_h_r_13')
// (10, 5, 'neigh_op_bnr_0')
// (11, 3, 'neigh_op_top_0')
// (11, 4, 'lutff_0/out')
// (11, 4, 'sp4_h_r_0')
// (11, 4, 'sp4_h_r_24')
// (11, 5, 'neigh_op_bot_0')
// (12, 3, 'neigh_op_tnl_0')
// (12, 4, 'neigh_op_lft_0')
// (12, 4, 'sp4_h_r_13')
// (12, 4, 'sp4_h_r_37')
// (12, 5, 'neigh_op_bnl_0')
// (13, 4, 'span4_horz_13')
// (13, 4, 'span4_horz_37')

reg n528 = 0;
// (9, 7, 'local_g0_0')
// (9, 7, 'lutff_6/in_0')
// (9, 7, 'sp4_h_r_8')
// (10, 6, 'neigh_op_tnr_0')
// (10, 7, 'neigh_op_rgt_0')
// (10, 7, 'sp4_h_r_21')
// (10, 8, 'neigh_op_bnr_0')
// (11, 6, 'local_g1_0')
// (11, 6, 'lutff_2/in_3')
// (11, 6, 'neigh_op_top_0')
// (11, 7, 'lutff_0/out')
// (11, 7, 'sp4_h_r_32')
// (11, 8, 'neigh_op_bot_0')
// (12, 6, 'neigh_op_tnl_0')
// (12, 7, 'neigh_op_lft_0')
// (12, 7, 'sp4_h_r_45')
// (12, 8, 'neigh_op_bnl_0')
// (13, 7, 'span4_horz_45')

reg n529 = 0;
// (9, 7, 'local_g0_2')
// (9, 7, 'lutff_2/in_0')
// (9, 7, 'sp4_h_r_10')
// (10, 6, 'neigh_op_tnr_1')
// (10, 7, 'neigh_op_rgt_1')
// (10, 7, 'sp4_h_r_23')
// (10, 8, 'neigh_op_bnr_1')
// (11, 6, 'neigh_op_top_1')
// (11, 7, 'lutff_1/out')
// (11, 7, 'sp4_h_r_34')
// (11, 8, 'neigh_op_bot_1')
// (12, 6, 'neigh_op_tnl_1')
// (12, 7, 'neigh_op_lft_1')
// (12, 7, 'sp4_h_r_47')
// (12, 8, 'neigh_op_bnl_1')
// (13, 7, 'span4_horz_47')

reg n530 = 0;
// (9, 9, 'local_g1_2')
// (9, 9, 'lutff_7/in_2')
// (9, 9, 'sp4_h_r_10')
// (10, 8, 'neigh_op_tnr_1')
// (10, 9, 'neigh_op_rgt_1')
// (10, 9, 'sp4_h_r_23')
// (10, 10, 'neigh_op_bnr_1')
// (11, 8, 'local_g1_1')
// (11, 8, 'lutff_7/in_3')
// (11, 8, 'neigh_op_top_1')
// (11, 9, 'local_g2_1')
// (11, 9, 'lutff_1/out')
// (11, 9, 'lutff_4/in_3')
// (11, 9, 'sp4_h_r_34')
// (11, 10, 'local_g0_1')
// (11, 10, 'lutff_4/in_1')
// (11, 10, 'neigh_op_bot_1')
// (12, 8, 'neigh_op_tnl_1')
// (12, 9, 'neigh_op_lft_1')
// (12, 9, 'sp4_h_r_47')
// (12, 10, 'neigh_op_bnl_1')
// (13, 9, 'span4_horz_47')

wire \d_out[1] ;
// (9, 10, 'sp4_h_r_0')
// (10, 9, 'neigh_op_tnr_4')
// (10, 10, 'neigh_op_rgt_4')
// (10, 10, 'sp4_h_r_13')
// (10, 11, 'neigh_op_bnr_4')
// (11, 9, 'neigh_op_top_4')
// (11, 10, 'lutff_4/out')
// (11, 10, 'sp4_h_r_24')
// (11, 11, 'neigh_op_bot_4')
// (12, 9, 'neigh_op_tnl_4')
// (12, 10, 'neigh_op_lft_4')
// (12, 10, 'sp4_h_r_37')
// (12, 11, 'neigh_op_bnl_4')
// (13, 10, 'span4_horz_37')
// (13, 10, 'span4_vert_t_14')
// (13, 11, 'span4_vert_b_14')
// (13, 12, 'io_0/D_OUT_0')
// (13, 12, 'io_0/PAD')
// (13, 12, 'local_g0_2')
// (13, 12, 'span4_vert_b_10')
// (13, 13, 'span4_vert_b_6')
// (13, 14, 'span4_vert_b_2')

reg n532 = 0;
// (9, 11, 'local_g1_0')
// (9, 11, 'lutff_7/in_0')
// (9, 11, 'sp4_h_r_8')
// (10, 10, 'neigh_op_tnr_0')
// (10, 11, 'neigh_op_rgt_0')
// (10, 11, 'sp4_h_r_21')
// (10, 12, 'neigh_op_bnr_0')
// (11, 10, 'neigh_op_top_0')
// (11, 11, 'lutff_0/out')
// (11, 11, 'sp4_h_r_32')
// (11, 12, 'neigh_op_bot_0')
// (12, 10, 'neigh_op_tnl_0')
// (12, 11, 'neigh_op_lft_0')
// (12, 11, 'sp4_h_r_45')
// (12, 12, 'neigh_op_bnl_0')
// (13, 11, 'span4_horz_45')

wire io_10_17_1;
// (9, 16, 'neigh_op_tnr_2')
// (9, 16, 'neigh_op_tnr_6')
// (10, 7, 'sp12_v_t_23')
// (10, 8, 'sp12_v_b_23')
// (10, 9, 'sp12_v_b_20')
// (10, 10, 'sp12_v_b_19')
// (10, 11, 'sp12_v_b_16')
// (10, 12, 'sp12_v_b_15')
// (10, 13, 'sp12_v_b_12')
// (10, 14, 'sp12_v_b_11')
// (10, 15, 'sp12_v_b_8')
// (10, 16, 'neigh_op_top_2')
// (10, 16, 'neigh_op_top_6')
// (10, 16, 'sp12_v_b_7')
// (10, 17, 'io_1/D_IN_0')
// (10, 17, 'io_1/PAD')
// (10, 17, 'span12_vert_4')
// (11, 16, 'neigh_op_tnl_2')
// (11, 16, 'neigh_op_tnl_6')

reg n534 = 0;
// (10, 2, 'neigh_op_tnr_2')
// (10, 3, 'neigh_op_rgt_2')
// (10, 4, 'neigh_op_bnr_2')
// (11, 2, 'neigh_op_top_2')
// (11, 3, 'local_g0_2')
// (11, 3, 'lutff_2/in_2')
// (11, 3, 'lutff_2/out')
// (11, 4, 'local_g0_2')
// (11, 4, 'local_g1_2')
// (11, 4, 'lutff_0/in_0')
// (11, 4, 'lutff_2/in_0')
// (11, 4, 'lutff_3/in_0')
// (11, 4, 'lutff_4/in_1')
// (11, 4, 'neigh_op_bot_2')
// (12, 2, 'neigh_op_tnl_2')
// (12, 3, 'neigh_op_lft_2')
// (12, 4, 'neigh_op_bnl_2')

reg n535 = 0;
// (10, 2, 'neigh_op_tnr_3')
// (10, 3, 'neigh_op_rgt_3')
// (10, 4, 'neigh_op_bnr_3')
// (11, 2, 'neigh_op_top_3')
// (11, 3, 'local_g0_3')
// (11, 3, 'lutff_3/in_2')
// (11, 3, 'lutff_3/out')
// (11, 4, 'local_g0_3')
// (11, 4, 'local_g1_3')
// (11, 4, 'lutff_0/in_1')
// (11, 4, 'lutff_2/in_1')
// (11, 4, 'lutff_3/in_1')
// (11, 4, 'lutff_4/in_0')
// (11, 4, 'neigh_op_bot_3')
// (12, 2, 'neigh_op_tnl_3')
// (12, 3, 'neigh_op_lft_3')
// (12, 4, 'neigh_op_bnl_3')

reg n536 = 0;
// (10, 2, 'neigh_op_tnr_4')
// (10, 2, 'sp4_r_v_b_37')
// (10, 3, 'neigh_op_rgt_4')
// (10, 3, 'sp4_r_v_b_24')
// (10, 4, 'neigh_op_bnr_4')
// (10, 4, 'sp4_r_v_b_13')
// (10, 5, 'sp4_r_v_b_0')
// (11, 1, 'sp4_v_t_37')
// (11, 2, 'neigh_op_top_4')
// (11, 2, 'sp4_v_b_37')
// (11, 3, 'local_g0_4')
// (11, 3, 'local_g1_4')
// (11, 3, 'lutff_1/in_2')
// (11, 3, 'lutff_4/in_2')
// (11, 3, 'lutff_4/out')
// (11, 3, 'sp4_v_b_24')
// (11, 4, 'local_g1_4')
// (11, 4, 'local_g1_5')
// (11, 4, 'lutff_0/in_2')
// (11, 4, 'lutff_2/in_2')
// (11, 4, 'lutff_3/in_2')
// (11, 4, 'lutff_4/in_2')
// (11, 4, 'neigh_op_bot_4')
// (11, 4, 'sp4_v_b_13')
// (11, 5, 'sp4_v_b_0')
// (12, 2, 'neigh_op_tnl_4')
// (12, 3, 'neigh_op_lft_4')
// (12, 4, 'neigh_op_bnl_4')

reg n537 = 0;
// (10, 2, 'neigh_op_tnr_7')
// (10, 3, 'neigh_op_rgt_7')
// (10, 4, 'neigh_op_bnr_7')
// (11, 2, 'neigh_op_top_7')
// (11, 3, 'local_g0_7')
// (11, 3, 'local_g1_7')
// (11, 3, 'lutff_0/in_1')
// (11, 3, 'lutff_4/in_3')
// (11, 3, 'lutff_7/in_3')
// (11, 3, 'lutff_7/out')
// (11, 4, 'local_g0_7')
// (11, 4, 'local_g1_7')
// (11, 4, 'lutff_0/in_3')
// (11, 4, 'lutff_2/in_3')
// (11, 4, 'lutff_3/in_3')
// (11, 4, 'lutff_4/in_3')
// (11, 4, 'neigh_op_bot_7')
// (12, 2, 'neigh_op_tnl_7')
// (12, 3, 'neigh_op_lft_7')
// (12, 4, 'neigh_op_bnl_7')

wire n538;
// (10, 3, 'neigh_op_tnr_1')
// (10, 4, 'neigh_op_rgt_1')
// (10, 5, 'neigh_op_bnr_1')
// (11, 2, 'sp4_r_v_b_43')
// (11, 3, 'local_g1_1')
// (11, 3, 'local_g1_6')
// (11, 3, 'lutff_2/in_0')
// (11, 3, 'lutff_3/in_0')
// (11, 3, 'lutff_4/in_0')
// (11, 3, 'neigh_op_top_1')
// (11, 3, 'sp4_r_v_b_30')
// (11, 4, 'lutff_1/out')
// (11, 4, 'sp4_r_v_b_19')
// (11, 5, 'neigh_op_bot_1')
// (11, 5, 'sp4_r_v_b_6')
// (12, 1, 'sp4_v_t_43')
// (12, 2, 'sp4_v_b_43')
// (12, 3, 'neigh_op_tnl_1')
// (12, 3, 'sp4_v_b_30')
// (12, 4, 'neigh_op_lft_1')
// (12, 4, 'sp4_v_b_19')
// (12, 5, 'neigh_op_bnl_1')
// (12, 5, 'sp4_v_b_6')

reg n539 = 0;
// (10, 4, 'neigh_op_tnr_0')
// (10, 5, 'neigh_op_rgt_0')
// (10, 6, 'neigh_op_bnr_0')
// (11, 4, 'neigh_op_top_0')
// (11, 5, 'local_g1_0')
// (11, 5, 'lutff_0/out')
// (11, 5, 'lutff_5/in_0')
// (11, 6, 'neigh_op_bot_0')
// (12, 4, 'neigh_op_tnl_0')
// (12, 5, 'neigh_op_lft_0')
// (12, 6, 'neigh_op_bnl_0')

reg n540 = 0;
// (10, 4, 'neigh_op_tnr_5')
// (10, 5, 'neigh_op_rgt_5')
// (10, 6, 'neigh_op_bnr_5')
// (11, 4, 'neigh_op_top_5')
// (11, 5, 'local_g1_5')
// (11, 5, 'lutff_2/in_0')
// (11, 5, 'lutff_5/out')
// (11, 6, 'neigh_op_bot_5')
// (12, 4, 'neigh_op_tnl_5')
// (12, 5, 'neigh_op_lft_5')
// (12, 6, 'neigh_op_bnl_5')

reg n541 = 0;
// (10, 5, 'neigh_op_tnr_6')
// (10, 6, 'neigh_op_rgt_6')
// (10, 7, 'neigh_op_bnr_6')
// (11, 5, 'neigh_op_top_6')
// (11, 6, 'local_g1_6')
// (11, 6, 'lutff_4/in_3')
// (11, 6, 'lutff_6/out')
// (11, 7, 'neigh_op_bot_6')
// (12, 5, 'neigh_op_tnl_6')
// (12, 6, 'neigh_op_lft_6')
// (12, 7, 'neigh_op_bnl_6')

reg n542 = 0;
// (10, 6, 'neigh_op_tnr_3')
// (10, 7, 'neigh_op_rgt_3')
// (10, 8, 'neigh_op_bnr_3')
// (11, 4, 'sp4_r_v_b_42')
// (11, 5, 'local_g1_7')
// (11, 5, 'lutff_0/in_0')
// (11, 5, 'sp4_r_v_b_31')
// (11, 6, 'neigh_op_top_3')
// (11, 6, 'sp4_r_v_b_18')
// (11, 7, 'lutff_3/out')
// (11, 7, 'sp4_r_v_b_7')
// (11, 8, 'neigh_op_bot_3')
// (12, 3, 'sp4_v_t_42')
// (12, 4, 'sp4_v_b_42')
// (12, 5, 'sp4_v_b_31')
// (12, 6, 'neigh_op_tnl_3')
// (12, 6, 'sp4_v_b_18')
// (12, 7, 'neigh_op_lft_3')
// (12, 7, 'sp4_v_b_7')
// (12, 8, 'neigh_op_bnl_3')

reg n543 = 0;
// (10, 6, 'neigh_op_tnr_7')
// (10, 7, 'neigh_op_rgt_7')
// (10, 8, 'neigh_op_bnr_7')
// (11, 6, 'neigh_op_top_7')
// (11, 7, 'local_g1_7')
// (11, 7, 'lutff_0/in_0')
// (11, 7, 'lutff_7/out')
// (11, 8, 'neigh_op_bot_7')
// (12, 6, 'neigh_op_tnl_7')
// (12, 7, 'neigh_op_lft_7')
// (12, 8, 'neigh_op_bnl_7')

reg n544 = 0;
// (10, 7, 'neigh_op_tnr_2')
// (10, 8, 'neigh_op_rgt_2')
// (10, 9, 'neigh_op_bnr_2')
// (11, 7, 'local_g1_2')
// (11, 7, 'lutff_7/in_0')
// (11, 7, 'neigh_op_top_2')
// (11, 8, 'lutff_2/out')
// (11, 9, 'neigh_op_bot_2')
// (12, 7, 'neigh_op_tnl_2')
// (12, 8, 'neigh_op_lft_2')
// (12, 9, 'neigh_op_bnl_2')

reg n545 = 0;
// (10, 7, 'neigh_op_tnr_7')
// (10, 8, 'neigh_op_rgt_7')
// (10, 9, 'neigh_op_bnr_7')
// (11, 7, 'local_g0_7')
// (11, 7, 'lutff_1/in_0')
// (11, 7, 'neigh_op_top_7')
// (11, 8, 'lutff_7/out')
// (11, 9, 'neigh_op_bot_7')
// (12, 7, 'neigh_op_tnl_7')
// (12, 8, 'neigh_op_lft_7')
// (12, 9, 'neigh_op_bnl_7')

reg n546 = 0;
// (10, 8, 'neigh_op_tnr_0')
// (10, 9, 'neigh_op_rgt_0')
// (10, 10, 'neigh_op_bnr_0')
// (11, 8, 'neigh_op_top_0')
// (11, 9, 'local_g1_0')
// (11, 9, 'lutff_0/out')
// (11, 9, 'lutff_1/in_0')
// (11, 10, 'neigh_op_bot_0')
// (12, 8, 'neigh_op_tnl_0')
// (12, 9, 'neigh_op_lft_0')
// (12, 10, 'neigh_op_bnl_0')

reg n547 = 0;
// (10, 8, 'neigh_op_tnr_4')
// (10, 9, 'neigh_op_rgt_4')
// (10, 10, 'neigh_op_bnr_4')
// (11, 8, 'neigh_op_top_4')
// (11, 9, 'lutff_4/out')
// (11, 10, 'local_g0_4')
// (11, 10, 'lutff_4/in_2')
// (11, 10, 'neigh_op_bot_4')
// (12, 8, 'neigh_op_tnl_4')
// (12, 9, 'neigh_op_lft_4')
// (12, 10, 'neigh_op_bnl_4')

reg n548 = 0;
// (10, 8, 'neigh_op_tnr_7')
// (10, 9, 'neigh_op_rgt_7')
// (10, 10, 'neigh_op_bnr_7')
// (11, 8, 'neigh_op_top_7')
// (11, 9, 'local_g1_7')
// (11, 9, 'lutff_0/in_0')
// (11, 9, 'lutff_7/out')
// (11, 10, 'neigh_op_bot_7')
// (12, 8, 'neigh_op_tnl_7')
// (12, 9, 'neigh_op_lft_7')
// (12, 10, 'neigh_op_bnl_7')

reg n549 = 0;
// (10, 10, 'neigh_op_tnr_1')
// (10, 11, 'neigh_op_rgt_1')
// (10, 12, 'neigh_op_bnr_1')
// (11, 10, 'neigh_op_top_1')
// (11, 11, 'local_g0_1')
// (11, 11, 'lutff_1/out')
// (11, 11, 'lutff_7/in_0')
// (11, 12, 'neigh_op_bot_1')
// (12, 10, 'neigh_op_tnl_1')
// (12, 11, 'neigh_op_lft_1')
// (12, 12, 'neigh_op_bnl_1')

reg n550 = 0;
// (10, 10, 'neigh_op_tnr_4')
// (10, 11, 'neigh_op_rgt_4')
// (10, 12, 'neigh_op_bnr_4')
// (11, 10, 'neigh_op_top_4')
// (11, 11, 'local_g0_4')
// (11, 11, 'lutff_0/in_0')
// (11, 11, 'lutff_4/out')
// (11, 12, 'neigh_op_bot_4')
// (12, 10, 'neigh_op_tnl_4')
// (12, 11, 'neigh_op_lft_4')
// (12, 12, 'neigh_op_bnl_4')

reg n551 = 0;
// (10, 10, 'neigh_op_tnr_5')
// (10, 11, 'neigh_op_rgt_5')
// (10, 12, 'neigh_op_bnr_5')
// (11, 10, 'neigh_op_top_5')
// (11, 11, 'local_g1_5')
// (11, 11, 'lutff_4/in_0')
// (11, 11, 'lutff_5/out')
// (11, 12, 'neigh_op_bot_5')
// (12, 10, 'neigh_op_tnl_5')
// (12, 11, 'neigh_op_lft_5')
// (12, 12, 'neigh_op_bnl_5')

reg n552 = 0;
// (10, 10, 'neigh_op_tnr_7')
// (10, 11, 'neigh_op_rgt_7')
// (10, 12, 'neigh_op_bnr_7')
// (11, 10, 'neigh_op_top_7')
// (11, 11, 'local_g1_7')
// (11, 11, 'lutff_5/in_3')
// (11, 11, 'lutff_7/out')
// (11, 12, 'neigh_op_bot_7')
// (12, 10, 'neigh_op_tnl_7')
// (12, 11, 'neigh_op_lft_7')
// (12, 12, 'neigh_op_bnl_7')

reg n553 = 0;
// (10, 11, 'neigh_op_tnr_7')
// (10, 12, 'neigh_op_rgt_7')
// (10, 13, 'neigh_op_bnr_7')
// (11, 11, 'local_g0_7')
// (11, 11, 'lutff_1/in_0')
// (11, 11, 'neigh_op_top_7')
// (11, 12, 'lutff_7/out')
// (11, 13, 'neigh_op_bot_7')
// (12, 11, 'neigh_op_tnl_7')
// (12, 12, 'neigh_op_lft_7')
// (12, 13, 'neigh_op_bnl_7')

wire n554;
// (11, 3, 'lutff_1/cout')
// (11, 3, 'lutff_2/in_3')

wire n555;
// (11, 3, 'lutff_2/cout')
// (11, 3, 'lutff_3/in_3')

wire n556;
// (2, 3, 'lutff_0/cout')

wire n557;
// (11, 3, 'lutff_0/cout')

wire n558;
// (5, 12, 'lutff_6/lout')

wire n559;
// (9, 12, 'lutff_1/lout')

wire n560;
// (2, 8, 'lutff_3/lout')

wire n561;
// (5, 4, 'lutff_2/lout')

wire n562;
// (6, 8, 'lutff_4/lout')

wire n563;
// (4, 8, 'lutff_5/lout')

wire n564;
// (7, 13, 'lutff_0/lout')

wire n565;
// (5, 5, 'lutff_3/lout')

wire n566;
// (2, 12, 'lutff_0/lout')

wire n567;
// (7, 5, 'lutff_5/lout')

wire n568;
// (6, 12, 'lutff_1/lout')

wire n569;
// (4, 12, 'lutff_2/lout')

wire n570;
// (9, 5, 'lutff_7/lout')

wire n571;
// (8, 15, 'lutff_5/lout')

wire n572;
// (5, 9, 'lutff_0/lout')

wire n573;
// (7, 9, 'lutff_2/lout')

wire n574;
// (9, 9, 'lutff_4/lout')

wire n575;
// (5, 8, 'lutff_4/lout')

wire n576;
// (7, 8, 'lutff_6/lout')

wire n577;
// (11, 3, 'lutff_3/lout')

wire n578;
// (6, 11, 'lutff_5/lout')

wire n579;
// (8, 11, 'lutff_7/lout')

wire n580;
// (5, 12, 'lutff_1/lout')

wire n581;
// (7, 1, 'lutff_3/lout')

wire n582;
// (4, 8, 'lutff_0/lout')

wire n583;
// (9, 12, 'lutff_5/lout')

wire n584;
// (2, 8, 'lutff_7/lout')

wire n585;
// (5, 4, 'lutff_6/lout')

wire n586;
// (7, 13, 'lutff_4/lout')

wire n587;
// (7, 5, 'lutff_0/lout')

wire n588;
// (9, 13, 'lutff_6/lout')

wire n589;
// (5, 5, 'lutff_7/lout')

wire n590;
// (4, 12, 'lutff_6/lout')

wire n591;
// (8, 4, 'lutff_3/lout')

wire n592;
// (8, 15, 'lutff_0/lout')

wire n593;
// (6, 7, 'lutff_3/lout')

wire n594;
// (8, 7, 'lutff_5/lout')

wire n595;
// (7, 8, 'lutff_1/lout')

wire n596;
// (9, 8, 'lutff_3/lout')

wire n597;
// (5, 11, 'lutff_4/lout')

wire n598;
// (4, 4, 'lutff_7/lout')

wire n599;
// (6, 11, 'lutff_0/lout')

wire n600;
// (8, 11, 'lutff_2/lout')

wire n601;
// (5, 12, 'lutff_5/lout')

wire n602;
// (6, 8, 'lutff_3/lout')

wire n603;
// (7, 1, 'lutff_7/lout')

wire n604;
// (4, 8, 'lutff_4/lout')

wire n605;
// (7, 12, 'lutff_7/lout')

wire n606;
// (6, 3, 'lutff_1/lout')

wire n607;
// (8, 3, 'lutff_3/lout')

wire n608;
// (1, 10, 'lutff_5/lout')

wire n609;
// (6, 6, 'lutff_6/lout')

wire n610;
// (8, 7, 'lutff_0/lout')

wire n611;
// (6, 7, 'lutff_7/lout')

wire n612;
// (5, 8, 'lutff_3/lout')

wire n613;
// (7, 8, 'lutff_5/lout')

wire n614;
// (6, 11, 'lutff_4/lout')

wire n615;
// (11, 6, 'lutff_4/lout')

wire n616;
// (11, 9, 'lutff_0/lout')

wire n617;
// (5, 12, 'lutff_0/lout')

wire n618;
// (7, 1, 'lutff_2/lout')

wire n619;
// (7, 12, 'lutff_2/lout')

wire n620;
// (9, 12, 'lutff_4/lout')

wire n621;
// (2, 11, 'lutff_2/lout')

wire n622;
// (6, 3, 'lutff_5/lout')

wire n623;
// (6, 6, 'lutff_1/lout')

wire n624;
// (8, 3, 'lutff_7/lout')

wire n625;
// (4, 11, 'lutff_0/lout')

wire n626;
// (9, 4, 'lutff_5/lout')

wire n627;
// (5, 7, 'lutff_6/lout')

wire n628;
// (9, 7, 'lutff_1/lout')

wire n629;
// (2, 3, 'lutff_3/lout')

wire n630;
// (4, 3, 'lutff_5/lout')

wire n631;
// (6, 7, 'lutff_2/lout')

wire n632;
// (8, 7, 'lutff_4/lout')

wire n633;
// (7, 8, 'lutff_0/lout')

wire n634;
// (5, 8, 'lutff_7/lout')

wire n635;
// (5, 11, 'lutff_3/lout')

wire n636;
// (7, 11, 'lutff_5/lout')

wire n637;
// (8, 11, 'lutff_1/lout')

wire n638;
// (6, 10, 'lutff_3/lout')

wire n639;
// (11, 9, 'lutff_4/lout')

wire n640;
// (8, 10, 'lutff_5/lout')

wire n641;
// (9, 11, 'lutff_3/lout')

wire n642;
// (5, 3, 'lutff_4/lout')

wire n643;
// (2, 10, 'lutff_1/lout')

wire n644;
// (7, 3, 'lutff_6/lout')

wire n645;
// (4, 10, 'lutff_3/lout')

wire n646;
// (6, 3, 'lutff_0/lout')

wire n647;
// (8, 3, 'lutff_2/lout')

wire n648;
// (8, 14, 'lutff_2/lout')

wire n649;
// (6, 6, 'lutff_5/lout')

wire n650;
// (9, 4, 'lutff_0/lout')

wire n651;
// (5, 7, 'lutff_1/lout')

wire n652;
// (4, 11, 'lutff_4/lout')

wire n653;
// (7, 7, 'lutff_3/lout')

wire n654;
// (2, 3, 'lutff_7/lout')

wire n655;
// (11, 5, 'lutff_2/lout')

wire n656;
// (5, 8, 'lutff_2/lout')

wire n657;
// (7, 8, 'lutff_4/lout')

wire n658;
// (9, 8, 'lutff_6/lout')

wire n659;
// (5, 11, 'lutff_7/lout')

wire n660;
// (4, 7, 'lutff_6/lout')

wire n661;
// (8, 10, 'lutff_0/lout')

wire n662;
// (6, 10, 'lutff_7/lout')

wire n663;
// (6, 2, 'lutff_3/lout')

wire n664;
// (8, 2, 'lutff_5/lout')

wire n665;
// (7, 3, 'lutff_1/lout')

wire n666;
// (9, 11, 'lutff_7/lout')

wire n667;
// (5, 6, 'lutff_4/lout')

wire n668;
// (4, 10, 'lutff_7/lout')

wire n669;
// (6, 3, 'lutff_4/lout')

wire n670;
// (6, 6, 'lutff_0/lout')

wire n671;
// (8, 3, 'lutff_6/lout')

wire n672;
// (8, 14, 'lutff_6/lout')

wire n673;
// (11, 4, 'lutff_5/lout')

wire n674;
// (9, 4, 'lutff_4/lout')

wire n675;
// (5, 7, 'lutff_5/lout')

wire n676;
// (9, 7, 'lutff_0/lout')

wire n677;
// (2, 14, 'lutff_2/lout')

wire n678;
// (7, 7, 'lutff_7/lout')

wire n679;
// (2, 3, 'lutff_2/lout')

wire n680;
// (6, 9, 'lutff_1/lout')

wire n681;
// (8, 6, 'lutff_7/lout')

wire n682;
// (2, 6, 'lutff_3/lout')

wire n683;
// (4, 6, 'lutff_5/lout')

wire n684;
// (6, 10, 'lutff_2/lout')

wire n685;
// (7, 14, 'lutff_6/lout')

wire n686;
// (8, 2, 'lutff_0/lout')

wire n687;
// (6, 2, 'lutff_7/lout')

wire n688;
// (6, 13, 'lutff_7/lout')

wire n689;
// (11, 8, 'lutff_7/lout')

wire n690;
// (5, 3, 'lutff_3/lout')

wire n691;
// (7, 3, 'lutff_5/lout')

wire n692;
// (4, 10, 'lutff_2/lout')

wire n693;
// (8, 3, 'lutff_1/lout')

wire n694;
// (6, 6, 'lutff_4/lout')

wire n695;
// (11, 4, 'lutff_0/lout')

wire n696;
// (5, 7, 'lutff_0/lout')

wire n697;
// (7, 7, 'lutff_2/lout')

wire n698;
// (5, 10, 'lutff_2/lout')

wire n699;
// (11, 5, 'lutff_1/lout')

wire n700;
// (8, 6, 'lutff_2/lout')

wire n701;
// (9, 10, 'lutff_6/lout')

wire n702;
// (5, 13, 'lutff_7/lout')

wire n703;
// (6, 9, 'lutff_5/lout')

wire n704;
// (4, 9, 'lutff_6/lout')

wire n705;
// (8, 9, 'lutff_7/lout')

wire n706;
// (6, 1, 'lutff_1/lout')

wire n707;
// (4, 6, 'lutff_0/lout')

wire n708;
// (5, 2, 'lutff_6/lout')

wire n709;
// (6, 10, 'lutff_6/lout')

wire n710;
// (6, 2, 'lutff_2/lout')

wire n711;
// (8, 2, 'lutff_4/lout')

wire n712;
// (11, 8, 'lutff_2/lout')

wire n713;
// (7, 3, 'lutff_0/lout')

wire n714;
// (9, 11, 'lutff_6/lout')

wire n715;
// (5, 3, 'lutff_7/lout')

wire n716;
// (5, 6, 'lutff_3/lout')

wire n717;
// (2, 2, 'lutff_0/lout')

wire n718;
// (6, 5, 'lutff_3/lout')

wire n719;
// (11, 4, 'lutff_4/lout')

wire n720;
// (8, 5, 'lutff_5/lout')

wire n721;
// (5, 10, 'lutff_6/lout')

wire n722;
// (5, 13, 'lutff_2/lout')

wire n723;
// (6, 9, 'lutff_0/lout')

wire n724;
// (8, 6, 'lutff_6/lout')

wire n725;
// (4, 9, 'lutff_1/lout')

wire n726;
// (8, 9, 'lutff_2/lout')

wire n727;
// (7, 2, 'lutff_4/lout')

wire n728;
// (5, 2, 'lutff_1/lout')

wire n729;
// (5, 14, 'lutff_3/lout')

wire n730;
// (4, 6, 'lutff_4/lout')

wire n731;
// (7, 14, 'lutff_5/lout')

wire n732;
// (6, 10, 'lutff_1/lout')

wire n733;
// (8, 10, 'lutff_3/lout')

wire n734;
// (6, 2, 'lutff_6/lout')

wire n735;
// (9, 11, 'lutff_1/lout')

wire n736;
// (5, 3, 'lutff_2/lout')

wire n737;
// (7, 3, 'lutff_4/lout')

wire n738;
// (5, 6, 'lutff_7/lout')

wire n739;
// (2, 2, 'lutff_4/lout')

wire n740;
// (7, 6, 'lutff_6/lout')

wire n741;
// (8, 13, 'lutff_4/lout')

wire n742;
// (8, 5, 'lutff_0/lout')

wire n743;
// (6, 5, 'lutff_7/lout')

wire n744;
// (11, 11, 'lutff_7/lout')

wire n745;
// (5, 10, 'lutff_1/lout')

wire n746;
// (8, 6, 'lutff_1/lout')

wire n747;
// (9, 10, 'lutff_5/lout')

wire n748;
// (5, 13, 'lutff_6/lout')

wire n749;
// (6, 9, 'lutff_4/lout')

wire n750;
// (4, 9, 'lutff_5/lout')

wire n751;
// (8, 9, 'lutff_6/lout')

wire n752;
// (11, 7, 'lutff_0/lout')

wire n753;
// (2, 6, 'lutff_6/lout')

wire n754;
// (5, 2, 'lutff_5/lout')

wire n755;
// (11, 8, 'lutff_1/lout')

wire n756;
// (1, 8, 'lutff_0/lout')

wire n757;
// (6, 12, 'lutff_5/lout')

wire n758;
// (7, 6, 'lutff_1/lout')

wire n759;
// (9, 6, 'lutff_3/lout')

wire n760;
// (5, 9, 'lutff_4/lout')

wire n761;
// (2, 5, 'lutff_1/lout')

wire n762;
// (6, 5, 'lutff_2/lout')

wire n763;
// (4, 5, 'lutff_3/lout')

wire n764;
// (8, 5, 'lutff_4/lout')

wire n765;
// (11, 3, 'lutff_7/lout')

wire n766;
// (5, 10, 'lutff_5/lout')

wire n767;
// (9, 10, 'lutff_0/lout')

wire n768;
// (7, 10, 'lutff_7/lout')

wire n769;
// (5, 13, 'lutff_1/lout')

wire n770;
// (7, 2, 'lutff_3/lout')

wire n771;
// (4, 9, 'lutff_0/lout')

wire n772;
// (8, 9, 'lutff_1/lout')

wire n773;
// (4, 6, 'lutff_3/lout')

wire n774;
// (9, 13, 'lutff_1/lout')

wire n775;
// (5, 5, 'lutff_2/lout')

wire n776;
// (7, 5, 'lutff_4/lout')

wire n777;
// (6, 12, 'lutff_0/lout')

wire n778;
// (4, 12, 'lutff_1/lout')

wire n779;
// (8, 4, 'lutff_7/lout')

wire n780;
// (7, 6, 'lutff_5/lout')

wire n781;
// (7, 9, 'lutff_1/lout')

wire n782;
// (8, 13, 'lutff_3/lout')

wire n783;
// (9, 9, 'lutff_3/lout')

wire n784;
// (6, 5, 'lutff_6/lout')

wire n785;
// (4, 5, 'lutff_7/lout')

wire n786;
// (11, 3, 'lutff_2/lout')

wire n787;
// (5, 10, 'lutff_0/lout')

wire n788;
// (7, 10, 'lutff_2/lout')

wire n789;
// (2, 9, 'lutff_2/lout')

wire n790;
// (7, 2, 'lutff_7/lout')

wire n791;
// (4, 9, 'lutff_4/lout')

wire n792;
// (6, 8, 'lutff_7/lout')

wire n793;
// (5, 5, 'lutff_6/lout')

wire n794;
// (9, 5, 'lutff_1/lout')

wire n795;
// (6, 12, 'lutff_4/lout')

wire n796;
// (6, 4, 'lutff_0/lout')

wire n797;
// (8, 4, 'lutff_2/lout')

wire n798;
// (7, 6, 'lutff_0/lout')

wire n799;
// (2, 13, 'lutff_4/lout')

wire n800;
// (5, 9, 'lutff_3/lout')

wire n801;
// (2, 5, 'lutff_0/lout')

wire n802;
// (7, 9, 'lutff_5/lout')

wire n803;
// (4, 13, 'lutff_6/lout')

wire n804;
// (4, 5, 'lutff_2/lout')

wire n805;
// (8, 5, 'lutff_3/lout')

wire n806;
// (9, 9, 'lutff_7/lout')

wire n807;
// (6, 5, 'lutff_1/lout')

wire n808;
// (11, 11, 'lutff_1/lout')

wire n809;
// (5, 12, 'lutff_4/lout')

wire n810;
// (7, 1, 'lutff_6/lout')

wire n811;
// (7, 12, 'lutff_6/lout')

wire n812;
// (4, 8, 'lutff_3/lout')

wire n813;
// (11, 7, 'lutff_3/lout')

wire n814;
// (11, 10, 'lutff_5/lout')

wire n815;
// (5, 5, 'lutff_1/lout')

wire n816;
// (7, 13, 'lutff_7/lout')

wire n817;
// (7, 5, 'lutff_3/lout')

wire n818;
// (9, 5, 'lutff_5/lout')

wire n819;
// (2, 4, 'lutff_3/lout')

wire n820;
// (6, 4, 'lutff_4/lout')

wire n821;
// (8, 4, 'lutff_6/lout')

wire n822;
// (6, 7, 'lutff_6/lout')

wire n823;
// (4, 13, 'lutff_1/lout')

wire n824;
// (7, 9, 'lutff_0/lout')

wire n825;
// (9, 6, 'lutff_6/lout')

wire n826;
// (9, 9, 'lutff_2/lout')

wire n827;
// (11, 11, 'lutff_5/lout')

wire n828;
// (11, 3, 'lutff_1/out')

wire n829;
// (11, 3, 'lutff_1/lout')

wire n830;
// (6, 11, 'lutff_3/lout')

wire n831;
// (8, 11, 'lutff_5/lout')

wire n832;
// (7, 1, 'lutff_1/lout')

wire n833;
// (7, 12, 'lutff_1/lout')

wire n834;
// (5, 4, 'lutff_4/lout')

wire n835;
// (6, 8, 'lutff_6/lout')

wire n836;
// (4, 8, 'lutff_7/lout')

wire n837;
// (7, 13, 'lutff_2/lout')

wire n838;
// (9, 13, 'lutff_4/lout')

wire n839;
// (5, 5, 'lutff_5/lout')

wire n840;
// (2, 12, 'lutff_2/lout')

wire n841;
// (7, 5, 'lutff_7/lout')

wire n842;
// (8, 4, 'lutff_1/lout')

wire n843;
// (2, 4, 'lutff_7/lout')

wire n844;
// (6, 7, 'lutff_1/lout')

wire n845;
// (8, 7, 'lutff_3/lout')

wire n846;
// (5, 8, 'lutff_6/lout')

wire n847;
// (5, 11, 'lutff_2/lout')

wire n848;
// (4, 4, 'lutff_5/lout')

wire n849;
// (8, 11, 'lutff_0/lout')

wire n850;
// (6, 11, 'lutff_7/lout')

wire n851;
// (11, 9, 'lutff_3/lout')

wire n852;
// (5, 12, 'lutff_3/lout')

wire n853;
// (2, 8, 'lutff_0/lout')

wire n854;
// (6, 8, 'lutff_1/lout')

wire n855;
// (7, 1, 'lutff_5/lout')

wire n856;
// (4, 8, 'lutff_2/lout')

wire n857;
// (7, 4, 'lutff_1/lout')

wire n858;
// (8, 8, 'lutff_3/lout')

wire n859;
// (7, 12, 'lutff_5/lout')

wire n860;
// (11, 10, 'lutff_4/lout')

wire n861;
// (5, 5, 'lutff_0/lout')

wire n862;
// (7, 5, 'lutff_2/lout')

wire n863;
// (4, 11, 'lutff_3/lout')

wire n864;
// (8, 15, 'lutff_2/lout')

wire n865;
// (2, 3, 'lutff_6/lout')

wire n866;
// (6, 7, 'lutff_5/lout')

wire n867;
// (8, 7, 'lutff_7/lout')

wire n868;
// (4, 4, 'lutff_0/lout')

wire n869;
// (5, 11, 'lutff_6/lout')

wire n870;
// (2, 7, 'lutff_3/lout')

wire n871;
// (6, 11, 'lutff_2/lout')

wire n872;
// (11, 6, 'lutff_2/lout')

wire n873;
// (8, 11, 'lutff_4/lout')

wire n874;
// (11, 9, 'lutff_7/lout')

wire n875;
// (7, 1, 'lutff_0/lout')

wire n876;
// (7, 12, 'lutff_0/lout')

wire n877;
// (5, 12, 'lutff_7/lout')

wire n878;
// (9, 12, 'lutff_2/lout')

wire n879;
// (4, 8, 'lutff_6/lout')

wire n880;
// (6, 3, 'lutff_3/lout')

wire n881;
// (8, 3, 'lutff_5/lout')

wire n882;
// (5, 7, 'lutff_4/lout')

wire n883;
// (2, 3, 'lutff_1/out')

wire n884;
// (2, 3, 'lutff_1/lout')

wire n885;
// (7, 7, 'lutff_6/lout')

wire n886;
// (4, 11, 'lutff_7/lout')

wire n887;
// (6, 7, 'lutff_0/lout')

wire n888;
// (8, 15, 'lutff_6/lout')

wire n889;
// (11, 5, 'lutff_5/lout')

wire n890;
// (7, 8, 'lutff_7/lout')

wire n891;
// (5, 11, 'lutff_1/lout')

wire n892;
// (11, 6, 'lutff_6/lout')

wire n893;
// (11, 9, 'lutff_2/lout')

wire n894;
// (7, 12, 'lutff_4/lout')

wire n895;
// (4, 8, 'lutff_1/lout')

wire n896;
// (7, 4, 'lutff_0/lout')

wire n897;
// (8, 3, 'lutff_0/lout')

wire n898;
// (8, 14, 'lutff_0/lout')

wire n899;
// (6, 3, 'lutff_7/lout')

wire n900;
// (6, 14, 'lutff_7/lout')

wire n901;
// (6, 6, 'lutff_3/lout')

wire n902;
// (9, 4, 'lutff_7/lout')

wire n903;
// (7, 7, 'lutff_1/lout')

wire n904;
// (9, 7, 'lutff_3/lout')

wire n905;
// (2, 3, 'lutff_5/lout')

wire n906;
// (4, 3, 'lutff_7/lout')

wire n907;
// (6, 7, 'lutff_4/lout')

wire n908;
// (8, 7, 'lutff_6/lout')

wire n909;
// (11, 13, 'lutff_4/lout')

wire n910;
// (11, 5, 'lutff_0/lout')

wire n911;
// (5, 8, 'lutff_0/lout')

wire n912;
// (7, 8, 'lutff_2/lout')

wire n913;
// (5, 11, 'lutff_5/lout')

wire n914;
// (7, 11, 'lutff_7/lout')

wire n915;
// (4, 7, 'lutff_4/lout')

wire n916;
// (6, 10, 'lutff_5/lout')

wire n917;
// (6, 2, 'lutff_1/lout')

wire n918;
// (6, 13, 'lutff_1/lout')

wire n919;
// (8, 10, 'lutff_7/lout')

wire n920;
// (8, 2, 'lutff_3/lout')

wire n921;
// (9, 11, 'lutff_5/lout')

wire n922;
// (5, 3, 'lutff_6/lout')

wire n923;
// (2, 10, 'lutff_3/lout')

wire n924;
// (5, 6, 'lutff_2/lout')

wire n925;
// (6, 3, 'lutff_2/lout')

wire n926;
// (8, 3, 'lutff_4/lout')

wire n927;
// (6, 6, 'lutff_7/lout')

wire n928;
// (11, 12, 'lutff_7/lout')

wire n929;
// (11, 4, 'lutff_3/lout')

wire n930;
// (9, 4, 'lutff_2/lout')

wire n931;
// (5, 7, 'lutff_3/lout')

wire n932;
// (2, 3, 'lutff_0/out')

wire n933;
// (2, 3, 'lutff_0/lout')

wire n934;
// (2, 3, 'carry_in_mux')

// Carry-In for (2 3)
assign n934 = 1;

wire n935;
// (4, 11, 'lutff_6/lout')

wire n936;
// (7, 7, 'lutff_5/lout')

wire n937;
// (4, 3, 'lutff_2/lout')

wire n938;
// (9, 7, 'lutff_7/lout')

wire n939;
// (8, 7, 'lutff_1/lout')

wire n940;
// (8, 6, 'lutff_5/lout')

wire n941;
// (5, 11, 'lutff_0/lout')

wire n942;
// (7, 11, 'lutff_2/lout')

wire n943;
// (5, 14, 'lutff_2/lout')

wire n944;
// (6, 10, 'lutff_0/lout')

wire n945;
// (11, 9, 'lutff_1/lout')

wire n946;
// (8, 10, 'lutff_2/lout')

wire n947;
// (6, 2, 'lutff_5/lout')

wire n948;
// (8, 2, 'lutff_7/lout')

wire n949;
// (9, 11, 'lutff_0/lout')

wire n950;
// (5, 3, 'lutff_1/lout')

wire n951;
// (7, 3, 'lutff_3/lout')

wire n952;
// (4, 10, 'lutff_0/lout')

wire n953;
// (9, 3, 'lutff_5/lout')

wire n954;
// (2, 10, 'lutff_7/lout')

wire n955;
// (5, 6, 'lutff_6/lout')

wire n956;
// (6, 3, 'lutff_6/lout')

wire n957;
// (6, 6, 'lutff_2/lout')

wire n958;
// (11, 12, 'lutff_2/lout')

wire n959;
// (11, 4, 'lutff_7/lout')

wire n960;
// (4, 11, 'lutff_1/lout')

wire n961;
// (7, 7, 'lutff_0/lout')

wire n962;
// (5, 7, 'lutff_7/lout')

wire n963;
// (9, 7, 'lutff_2/lout')

wire n964;
// (2, 3, 'lutff_4/lout')

wire n965;
// (2, 14, 'lutff_4/lout')

wire n966;
// (4, 14, 'lutff_6/lout')

wire n967;
// (8, 6, 'lutff_0/lout')

wire n968;
// (6, 9, 'lutff_3/lout')

wire n969;
// (8, 9, 'lutff_5/lout')

wire n970;
// (5, 2, 'lutff_4/lout')

wire n971;
// (5, 14, 'lutff_6/lout')

wire n972;
// (4, 6, 'lutff_7/lout')

wire n973;
// (6, 10, 'lutff_4/lout')

wire n974;
// (6, 2, 'lutff_0/lout')

wire n975;
// (8, 10, 'lutff_6/lout')

wire n976;
// (8, 2, 'lutff_2/lout')

wire n977;
// (9, 11, 'lutff_4/lout')

wire n978;
// (5, 3, 'lutff_5/lout')

wire n979;
// (7, 3, 'lutff_7/lout')

wire n980;
// (5, 6, 'lutff_1/lout')

wire n981;
// (4, 2, 'lutff_0/lout')

wire n982;
// (8, 13, 'lutff_7/lout')

wire n983;
// (11, 4, 'lutff_2/lout')

wire n984;
// (9, 4, 'lutff_1/lout')

wire n985;
// (1, 12, 'lutff_5/lout')

wire n986;
// (5, 7, 'lutff_2/lout')

wire n987;
// (7, 7, 'lutff_4/lout')

wire n988;
// (4, 3, 'lutff_1/lout')

wire n989;
// (4, 14, 'lutff_1/lout')

wire n990;
// (9, 7, 'lutff_6/lout')

wire n991;
// (5, 10, 'lutff_4/lout')

wire n992;
// (5, 13, 'lutff_0/lout')

wire n993;
// (8, 6, 'lutff_4/lout')

wire n994;
// (7, 2, 'lutff_2/lout')

wire n995;
// (8, 9, 'lutff_0/lout')

wire n996;
// (6, 9, 'lutff_7/lout')

wire n997;
// (4, 6, 'lutff_2/lout')

wire n998;
// (8, 10, 'lutff_1/lout')

wire n999;
// (6, 2, 'lutff_4/lout')

wire n1000;
// (6, 13, 'lutff_4/lout')

wire n1001;
// (8, 2, 'lutff_6/lout')

wire n1002;
// (5, 3, 'lutff_0/lout')

wire n1003;
// (7, 3, 'lutff_2/lout')

wire n1004;
// (5, 6, 'lutff_5/lout')

wire n1005;
// (7, 6, 'lutff_4/lout')

wire n1006;
// (8, 13, 'lutff_2/lout')

wire n1007;
// (6, 5, 'lutff_5/lout')

wire n1008;
// (11, 4, 'lutff_6/lout')

wire n1009;
// (8, 5, 'lutff_7/lout')

wire n1010;
// (9, 10, 'lutff_3/lout')

wire n1011;
// (5, 13, 'lutff_4/lout')

wire n1012;
// (6, 9, 'lutff_2/lout')

wire n1013;
// (7, 2, 'lutff_6/lout')

wire n1014;
// (4, 9, 'lutff_3/lout')

wire n1015;
// (8, 9, 'lutff_4/lout')

wire n1016;
// (11, 7, 'lutff_7/lout')

wire n1017;
// (5, 2, 'lutff_3/lout')

wire n1018;
// (5, 14, 'lutff_5/lout')

wire n1019;
// (7, 14, 'lutff_7/lout')

wire n1020;
// (8, 2, 'lutff_1/lout')

wire n1021;
// (6, 12, 'lutff_3/lout')

wire n1022;
// (8, 12, 'lutff_5/lout')

wire n1023;
// (5, 6, 'lutff_0/lout')

wire n1024;
// (9, 6, 'lutff_1/lout')

wire n1025;
// (5, 9, 'lutff_2/lout')

wire n1026;
// (4, 13, 'lutff_5/lout')

wire n1027;
// (8, 13, 'lutff_6/lout')

wire n1028;
// (6, 5, 'lutff_0/lout')

wire n1029;
// (11, 4, 'lutff_1/lout')

wire n1030;
// (7, 9, 'lutff_4/lout')

wire n1031;
// (8, 5, 'lutff_2/lout')

wire n1032;
// (9, 9, 'lutff_6/lout')

wire n1033;
// (11, 11, 'lutff_0/lout')

wire n1034;
// (5, 10, 'lutff_3/lout')

wire n1035;
// (7, 10, 'lutff_5/lout')

wire n1036;
// (8, 6, 'lutff_3/lout')

wire n1037;
// (7, 2, 'lutff_1/lout')

wire n1038;
// (9, 10, 'lutff_7/lout')

wire n1039;
// (2, 9, 'lutff_5/lout')

wire n1040;
// (6, 9, 'lutff_6/lout')

wire n1041;
// (4, 9, 'lutff_7/lout')

wire n1042;
// (4, 6, 'lutff_1/lout')

wire n1043;
// (7, 14, 'lutff_2/lout')

wire n1044;
// (5, 2, 'lutff_7/lout')

wire n1045;
// (7, 13, 'lutff_6/lout')

wire n1046;
// (8, 12, 'lutff_0/lout')

wire n1047;
// (1, 8, 'lutff_2/lout')

wire n1048;
// (6, 12, 'lutff_7/lout')

wire n1049;
// (6, 4, 'lutff_3/lout')

wire n1050;
// (8, 4, 'lutff_5/lout')

wire n1051;
// (7, 6, 'lutff_3/lout')

wire n1052;
// (8, 13, 'lutff_1/lout')

wire n1053;
// (9, 6, 'lutff_5/lout')

wire n1054;
// (5, 9, 'lutff_6/lout')

wire n1055;
// (9, 9, 'lutff_1/lout')

wire n1056;
// (2, 5, 'lutff_3/lout')

wire n1057;
// (6, 5, 'lutff_4/lout')

wire n1058;
// (4, 5, 'lutff_5/lout')

wire n1059;
// (8, 5, 'lutff_6/lout')

wire n1060;
// (11, 11, 'lutff_4/lout')

wire n1061;
// (11, 3, 'lutff_0/out')

wire n1062;
// (11, 3, 'lutff_0/lout')

wire n1063;
// (11, 3, 'carry_in_mux')

// Carry-In for (11 3)
assign n1063 = 1;

wire n1064;
// (7, 10, 'lutff_0/lout')

wire n1065;
// (5, 10, 'lutff_7/lout')

wire n1066;
// (9, 10, 'lutff_2/lout')

wire n1067;
// (7, 2, 'lutff_5/lout')

wire n1068;
// (4, 9, 'lutff_2/lout')

wire n1069;
// (8, 9, 'lutff_3/lout')

wire n1070;
// (5, 2, 'lutff_2/lout')

wire n1071;
// (7, 13, 'lutff_1/lout')

wire n1072;
// (5, 5, 'lutff_4/lout')

wire n1073;
// (7, 5, 'lutff_6/lout')

wire n1074;
// (6, 12, 'lutff_2/lout')

wire n1075;
// (4, 12, 'lutff_3/lout')

wire n1076;
// (8, 4, 'lutff_0/lout')

wire n1077;
// (2, 4, 'lutff_6/lout')

wire n1078;
// (6, 4, 'lutff_7/lout')

wire n1079;
// (9, 6, 'lutff_0/lout')

wire n1080;
// (5, 9, 'lutff_1/lout')

wire n1081;
// (7, 6, 'lutff_7/lout')

wire n1082;
// (8, 13, 'lutff_5/lout')

wire n1083;
// (7, 9, 'lutff_3/lout')

wire n1084;
// (4, 5, 'lutff_0/lout')

wire n1085;
// (8, 5, 'lutff_1/lout')

wire n1086;
// (9, 9, 'lutff_5/lout')

wire n1087;
// (11, 3, 'lutff_4/lout')

wire n1088;
// (7, 2, 'lutff_0/lout')

wire n1089;
// (7, 1, 'lutff_4/lout')

wire n1090;
// (11, 7, 'lutff_1/lout')

wire n1091;
// (5, 4, 'lutff_7/lout')

wire n1092;
// (7, 13, 'lutff_5/lout')

wire n1093;
// (7, 5, 'lutff_1/lout')

wire n1094;
// (2, 12, 'lutff_5/lout')

wire n1095;
// (6, 12, 'lutff_6/lout')

wire n1096;
// (2, 4, 'lutff_1/lout')

wire n1097;
// (4, 12, 'lutff_7/lout')

wire n1098;
// (6, 4, 'lutff_2/lout')

wire n1099;
// (8, 4, 'lutff_4/lout')

wire n1100;
// (11, 2, 'lutff_7/lout')

wire n1101;
// (7, 6, 'lutff_2/lout')

wire n1102;
// (9, 6, 'lutff_4/lout')

wire n1103;
// (5, 9, 'lutff_5/lout')

wire n1104;
// (9, 9, 'lutff_0/lout')

wire n1105;
// (2, 5, 'lutff_2/lout')

wire n1106;
// (7, 9, 'lutff_7/lout')

wire n1107;
// (4, 5, 'lutff_4/lout')

wire n1108;
// (11, 11, 'lutff_3/lout')

wire n1109;
// (6, 11, 'lutff_1/lout')

wire n1110;
// (8, 11, 'lutff_3/lout')

assign n829  = /* LUT   11  3  1 */ 1'b0;
assign n884  = /* LUT    2  3  1 */ 1'b0;
assign n933  = /* LUT    2  3  0 */ 1'b0;
assign n1062 = /* LUT   11  3  0 */ 1'b0;
assign n558  = /* LUT    5 12  6 */ n226;
assign n559  = /* LUT    9 12  1 */ n324;
assign n560  = /* LUT    2  8  3 */ (n19 ? n33 : n70);
assign n561  = /* LUT    5  4  2 */ n166;
assign n562  = /* LUT    6  8  4 */ n295;
assign n563  = /* LUT    4  8  5 */ (n170 ? (n46 ? n75 : 1'b0) : (n46 ? !n75 : 1'b1));
assign n564  = /* LUT    7 13  0 */ (n18 ? (n15 ? 1'b1 : !n398) : (n15 ? !n402 : 1'b1));
assign n565  = /* LUT    5  5  3 */ (n175 ? (n263 ? (n169 ? !n258 : 1'b1) : (n169 ? n258 : 1'b0)) : (n263 ? (n169 ? n258 : 1'b0) : (n169 ? !n258 : 1'b1)));
assign n566  = /* LUT    2 12  0 */ (n15 ? (n18 ? n82 : n98) : n82);
assign n567  = /* LUT    7  5  5 */ (n361 ? (n274 ? (n270 ? !n269 : 1'b0) : (n270 ? 1'b0 : !n269)) : (n274 ? (n270 ? n269 : 1'b0) : (n270 ? 1'b0 : n269)));
assign n568  = /* LUT    6 12  1 */ n304;
assign n569  = /* LUT    4 12  2 */ n50;
assign n570  = /* LUT    9  5  7 */ n350;
assign n571  = /* LUT    8 15  5 */ n478;
assign n572  = /* LUT    5  9  0 */ (n192 ? (n221 ? (n293 ? !n39 : 1'b1) : (n293 ? 1'b1 : !n39)) : 1'b0);
assign n573  = /* LUT    7  9  2 */ n380;
assign n574  = /* LUT    9  9  4 */ n507;
assign n575  = /* LUT    5  8  4 */ (n174 ? !n183 : n183);
assign n576  = /* LUT    7  8  6 */ (n188 ? (n46 ? !n371 : 1'b1) : (n46 ? n371 : 1'b0));
assign n577  = /* LUT   11  3  3 */ (n555 ? (n535 ? 1'b0 : !n538) : (n535 ? !n538 : 1'b0));
assign n578  = /* LUT    6 11  5 */ (n174 ? (n178 ? (n308 ? !n46 : 1'b1) : (n308 ? n46 : 1'b0)) : (n178 ? (n308 ? n46 : 1'b0) : (n308 ? !n46 : 1'b1)));
assign n579  = /* LUT    8 11  7 */ n465;
assign n580  = /* LUT    5 12  1 */ (n222 ? (n18 ? (n15 ? !n53 : 1'b1) : 1'b1) : 1'b0);
assign n581  = /* LUT    7  1  3 */ (n407 ? (n336 ? 1'b0 : (n334 ? n328 : 1'b1)) : 1'b0);
assign n582  = /* LUT    4  8  0 */ (n19 ? !n125 : !n34);
assign n583  = /* LUT    9 12  5 */ n522;
assign n584  = /* LUT    2  8  7 */ (n19 ? n75 : n26);
assign n585  = /* LUT    5  4  6 */ (n240 ? (n157 ? n14 : 1'b1) : (n157 ? !n14 : 1'b0));
assign n586  = /* LUT    7 13  4 */ n401;
assign n587  = /* LUT    7  5  0 */ (n363 ? (n357 ? (n274 ? n361 : 1'b1) : (n274 ? !n361 : 1'b0)) : (n357 ? (n274 ? !n361 : 1'b0) : (n274 ? n361 : 1'b1)));
assign n588  = /* LUT    9 13  6 */ n524;
assign n589  = /* LUT    5  5  7 */ (n17 ? !n67 : n67);
assign n590  = /* LUT    4 12  6 */ (n18 ? (n15 ? n142 : n98) : n142);
assign n591  = /* LUT    8  4  3 */ (n423 ? (n422 ? (n420 ? !n431 : n431) : (n420 ? n431 : !n431)) : (n422 ? (n420 ? n431 : !n431) : (n420 ? !n431 : n431)));
assign n592  = /* LUT    8 15  0 */ n483;
assign n593  = /* LUT    6  7  3 */ (n133 ? (n136 ? n149 : !n149) : (n136 ? !n149 : n149));
assign n594  = /* LUT    8  7  5 */ (n443 ? !n40 : !n450);
assign n595  = /* LUT    7  8  1 */ (n19 ? n373 : n288);
assign n596  = /* LUT    9  8  3 */ (n32 ? !n268 : n268);
assign n597  = /* LUT    5 11  4 */ (n19 ? n215 : n220);
assign n598  = /* LUT    4  4  7 */ n114;
assign n599  = /* LUT    6 11  0 */ (n19 ? !n311 : !n313);
assign n600  = /* LUT    8 11  2 */ (n481 ? (n48 ? n14 : 1'b1) : (n48 ? !n14 : 1'b0));
assign n601  = /* LUT    5 12  5 */ (n39 ? n51 : (n96 ? n214 : !n214));
assign n602  = /* LUT    6  8  3 */ (n285 ? (n378 ? (n30 ? !n39 : 1'b1) : (n30 ? 1'b1 : !n39)) : 1'b0);
assign n603  = /* LUT    7  1  7 */ (n340 ? (n327 ? !n338 : n338) : (n327 ? n338 : !n338));
assign n604  = /* LUT    4  8  4 */ (n193 ? (n46 ? !n33 : 1'b1) : (n46 ? n33 : 1'b0));
assign n605  = /* LUT    7 12  7 */ n389;
assign n606  = /* LUT    6  3  1 */ (n253 ? !n347 : n347);
assign n607  = /* LUT    8  3  3 */ (n427 ? 1'b0 : !n424);
assign n608  = /* LUT    1 10  5 */ n78;
assign n609  = /* LUT    6  6  6 */ (n279 ? (n169 ? (n68 ? n272 : !n272) : (n68 ? !n272 : n272)) : (n169 ? (n68 ? !n272 : n272) : (n68 ? n272 : !n272)));
assign n610  = /* LUT    8  7  0 */ (n13 ? 1'b0 : (n283 ? 1'b0 : !n419));
assign n611  = /* LUT    6  7  7 */ (n39 ? n199 : (n29 ? n292 : !n292));
assign n612  = /* LUT    5  8  3 */ (n172 ? !n170 : n170);
assign n613  = /* LUT    7  8  5 */ (n32 ? (n46 ? !n373 : 1'b1) : (n46 ? n373 : 1'b0));
assign n614  = /* LUT    6 11  4 */ (n178 ? (n46 ? n309 : 1'b0) : (n46 ? !n309 : 1'b1));
assign n615  = /* LUT   11  6  4 */ (n541 ? (n13 ? 1'b1 : (n283 ? 1'b1 : n419)) : 1'b0);
assign n616  = /* LUT   11  9  0 */ n548;
assign n617  = /* LUT    5 12  0 */ (n18 ? (n15 ? 1'b1 : !n235) : (n15 ? !n218 : 1'b1));
assign n618  = /* LUT    7  1  2 */ (n340 ? (n327 ? (n338 ? !n84 : 1'b0) : (n338 ? 1'b0 : !n84)) : (n327 ? (n338 ? 1'b0 : !n84) : (n338 ? !n84 : 1'b0)));
assign n619  = /* LUT    7 12  2 */ n385;
assign n620  = /* LUT    9 12  4 */ n96;
assign n621  = /* LUT    2 11  2 */ n45;
assign n622  = /* LUT    6  3  5 */ (n256 ? !n348 : n348);
assign n623  = /* LUT    6  6  1 */ (n149 ? (n276 ? n273 : !n273) : (n276 ? !n273 : n273));
assign n624  = /* LUT    8  3  7 */ (n420 ? !n432 : n432);
assign n625  = /* LUT    4 11  0 */ (n18 ? (n15 ? 1'b1 : !n142) : (n15 ? !n82 : 1'b1));
assign n626  = /* LUT    9  4  5 */ (rst ? 1'b0 : (n283 ? 1'b1 : (n13 ? !n434 : 1'b0)));
assign n627  = /* LUT    5  7  6 */ n197;
assign n628  = /* LUT    9  7  1 */ n497;
assign n629  = /* LUT    2  3  3 */ (n86 ? !n58 : n58);
assign n630  = /* LUT    4  3  5 */ (n59 ? !n11 : 1'b0);
assign n631  = /* LUT    6  7  2 */ (n280 ? (n29 ? (n292 ? !n39 : 1'b1) : (n292 ? 1'b1 : !n39)) : 1'b0);
assign n632  = /* LUT    8  7  4 */ (n198 ? (n13 ? 1'b0 : (n283 ? 1'b0 : !n419)) : 1'b0);
assign n633  = /* LUT    7  8  0 */ (n32 ? (n46 ? !n375 : 1'b1) : (n46 ? n375 : 1'b0));
assign n634  = /* LUT    5  8  7 */ n204;
assign n635  = /* LUT    5 11  3 */ (n200 ? (n45 ? n46 : 1'b0) : (n45 ? !n46 : 1'b1));
assign n636  = /* LUT    7 11  5 */ (n395 ? !n349 : n349);
assign n637  = /* LUT    8 11  1 */ n468;
assign n638  = /* LUT    6 10  3 */ (n174 ? (n46 ? !n301 : 1'b1) : (n46 ? n301 : 1'b0));
assign n639  = /* LUT   11  9  4 */ (n530 ? (n188 ? n250 : !n250) : (n188 ? !n250 : n250));
assign n640  = /* LUT    8 10  5 */ n460;
assign n641  = /* LUT    9 11  3 */ n464;
assign n642  = /* LUT    5  3  4 */ (n92 ? (n103 ? !n252 : n252) : 1'b0);
assign n643  = /* LUT    2 10  1 */ n35;
assign n644  = /* LUT    7  3  6 */ (n418 ? (n413 ? 1'b1 : n330) : (n413 ? n242 : (n330 ? n242 : !n242)));
assign n645  = /* LUT    4 10  3 */ (n19 ? !n127 : !n132);
assign n646  = /* LUT    6  3  0 */ (n92 ? (n154 ? (n255 ? !n254 : n254) : (n255 ? n254 : !n254)) : 1'b0);
assign n647  = /* LUT    8  3  2 */ (n430 ? !n432 : n432);
assign n648  = /* LUT    8 14  2 */ n479;
assign n649  = /* LUT    6  6  5 */ (n136 ? (n149 ? n278 : !n278) : (n149 ? !n278 : n278));
assign n650  = /* LUT    9  4  0 */ (n13 ? (n434 ? (n488 ? n527 : 1'b1) : 1'b0) : (n488 ? n527 : 1'b1));
assign n651  = /* LUT    5  7  1 */ (n23 ? (n181 ? n183 : !n183) : (n181 ? !n183 : n183));
assign n652  = /* LUT    4 11  4 */ n141;
assign n653  = /* LUT    7  7  3 */ n370;
assign n654  = /* LUT    2  3  7 */ (n90 ? !n11 : n11);
assign n655  = /* LUT   11  5  2 */ n540;
assign n656  = /* LUT    5  8  2 */ (n178 ? (n172 ? !n170 : n170) : (n172 ? n170 : !n170));
assign n657  = /* LUT    7  8  4 */ (n19 ? n375 : n372);
assign n658  = /* LUT    9  8  6 */ n29;
assign n659  = /* LUT    5 11  7 */ (n19 ? n216 : n49);
assign n660  = /* LUT    4  7  6 */ n121;
assign n661  = /* LUT    8 10  0 */ n457;
assign n662  = /* LUT    6 10  7 */ (n170 ? (n46 ? n302 : 1'b0) : (n46 ? !n302 : 1'b1));
assign n663  = /* LUT    6  2  3 */ (n333 ? (n84 ? (n334 ? 1'b1 : n335) : (n334 ? n335 : 1'b1)) : (n84 ? 1'b0 : n335));
assign n664  = /* LUT    8  2  5 */ (n421 ? n415 : !n415);
assign n665  = /* LUT    7  3  1 */ (n8 ? (n339 ? !n243 : n243) : (n339 ? n243 : !n243));
assign n666  = /* LUT    9 11  7 */ n532;
assign n667  = /* LUT    5  6  4 */ (n68 ? (n94 ? (n275 ? !n259 : n259) : n259) : (n94 ? n275 : 1'b1));
assign n668  = /* LUT    4 10  7 */ (n138 ? (n24 ? (n134 ? !n39 : 1'b1) : (n134 ? 1'b1 : !n39)) : 1'b0);
assign n669  = /* LUT    6  3  4 */ (n12 ? n251 : !n251);
assign n670  = /* LUT    6  6  0 */ (n169 ? n68 : !n68);
assign n671  = /* LUT    8  3  6 */ (n414 ? (n417 ? n91 : !n91) : (n417 ? !n91 : n91));
assign n672  = /* LUT    8 14  6 */ n480;
assign n673  = /* LUT   11  4  5 */ (n13 ? 1'b0 : !n419);
assign n674  = /* LUT    9  4  4 */ (rst ? 1'b0 : (n5 ? 1'b1 : (n488 ? !n527 : 1'b0)));
assign n675  = /* LUT    5  7  5 */ n196;
assign n676  = /* LUT    9  7  0 */ n498;
assign n677  = /* LUT    2 14  2 */ n54;
assign n678  = /* LUT    7  7  7 */ n198;
assign n679  = /* LUT    2  3  2 */ (n85 ? !n57 : n57);
assign n680  = /* LUT    6  9  1 */ (n19 ? !n299 : !n294);
assign n681  = /* LUT    8  6  7 */ n38;
assign n682  = /* LUT    2  6  3 */ n25;
assign n683  = /* LUT    4  6  5 */ !n65;
assign n684  = /* LUT    6 10  2 */ (n174 ? (n46 ? !n303 : 1'b1) : (n46 ? n303 : 1'b0));
assign n685  = /* LUT    7 14  6 */ n403;
assign n686  = /* LUT    8  2  0 */ (n410 ? (n162 ? (n341 ? 1'b0 : n407) : (n341 ? n407 : 1'b0)) : (n162 ? (n341 ? 1'b1 : !n407) : (n341 ? !n407 : 1'b1)));
assign n687  = /* LUT    6  2  7 */ (n342 ? (n239 ? n249 : 1'b1) : (n239 ? (n249 ? !n244 : n244) : n244));
assign n688  = /* LUT    6 13  7 */ n322;
assign n689  = /* LUT   11  8  7 */ (n530 ? !n250 : n250);
assign n690  = /* LUT    5  3  3 */ (n159 ? (n59 ? (n11 ? 1'b0 : !n9) : n11) : 1'b0);
assign n691  = /* LUT    7  3  5 */ (n108 ? (n417 ? n330 : 1'b1) : (n417 ? (n330 ? n242 : !n242) : n242));
assign n692  = /* LUT    4 10  2 */ (n19 ? !n131 : !n130);
assign n693  = /* LUT    8  3  1 */ (n421 ? !n249 : n249);
assign n694  = /* LUT    6  6  4 */ (n149 ? (n278 ? !n286 : n286) : (n278 ? n286 : !n286));
assign n695  = /* LUT   11  4  0 */ (n537 ? (n536 ? 1'b0 : (n535 ? 1'b0 : !n534)) : 1'b0);
assign n696  = /* LUT    5  7  0 */ (n23 ? n171 : !n171);
assign n697  = /* LUT    7  7  2 */ n120;
assign n698  = /* LUT    5 10  2 */ n208;
assign n699  = /* LUT   11  5  1 */ (rst ? 1'b1 : (n66 ? !n185 : 1'b0));
assign n700  = /* LUT    8  6  2 */ (n495 ? (n13 ? 1'b0 : (n283 ? 1'b0 : !n419)) : 1'b0);
assign n701  = /* LUT    9 10  6 */ n513;
assign n702  = /* LUT    5 13  7 */ n232;
assign n703  = /* LUT    6  9  5 */ (n200 ? (n188 ? (n295 ? !n46 : 1'b1) : (n295 ? n46 : 1'b0)) : (n188 ? (n295 ? n46 : 1'b0) : (n295 ? !n46 : 1'b1)));
assign n704  = /* LUT    4  9  6 */ (n19 ? n124 : n71);
assign n705  = /* LUT    8  9  7 */ (n15 ? (n18 ? n454 : n461) : n454);
assign n706  = /* LUT    6  1  1 */ (n335 ? n328 : (n333 ? 1'b1 : n334));
assign n707  = /* LUT    4  6  0 */ (n178 ? n25 : !n25);
assign n708  = /* LUT    5  2  6 */ (n241 ? (n151 ? !n7 : 1'b1) : (n151 ? n7 : 1'b0));
assign n709  = /* LUT    6 10  6 */ (n19 ? n303 : n305);
assign n710  = /* LUT    6  2  2 */ (n248 ? (n344 ? (n12 ? !n246 : n246) : (n12 ? n246 : !n246)) : (n344 ? (n12 ? n246 : !n246) : (n12 ? !n246 : n246)));
assign n711  = /* LUT    8  2  4 */ (n412 ? n340 : !n340);
assign n712  = /* LUT   11  8  2 */ n345;
assign n713  = /* LUT    7  3  0 */ (n343 ? (n105 ? (n251 ? 1'b1 : !n92) : (n251 ? !n92 : 1'b1)) : (n105 ? (n251 ? 1'b0 : n92) : (n251 ? n92 : 1'b0)));
assign n714  = /* LUT    9 11  6 */ n466;
assign n715  = /* LUT    5  3  7 */ (n170 ? n157 : !n157);
assign n716  = /* LUT    5  6  3 */ (n122 ? (n179 ? n123 : !n123) : (n179 ? !n123 : n123));
assign n717  = /* LUT    2  2  0 */ (n9 ? (n11 ? n7 : 1'b0) : 1'b0);
assign n718  = /* LUT    6  5  3 */ (n361 ? (n269 ? 1'b1 : n264) : (n269 ? n267 : (n264 ? n267 : !n267)));
assign n719  = /* LUT   11  4  4 */ (n537 ? (n536 ? (n534 ? !n535 : 1'b0) : 1'b0) : 1'b0);
assign n720  = /* LUT    8  5  5 */ (n444 ? 1'b0 : !n446);
assign n721  = /* LUT    5 10  6 */ n207;
assign n722  = /* LUT    5 13  2 */ (n15 ? (n18 ? n231 : n51) : n231);
assign n723  = /* LUT    6  9  0 */ (n18 ? (n15 ? 1'b1 : !n320) : (n15 ? !n41 : 1'b1));
assign n724  = /* LUT    8  6  6 */ n24;
assign n725  = /* LUT    4  9  1 */ (n193 ? (n46 ? !n124 : 1'b1) : (n46 ? n124 : 1'b0));
assign n726  = /* LUT    8  9  2 */ (n18 ? (n15 ? 1'b1 : !n451) : (n15 ? !n454 : 1'b1));
assign n727  = /* LUT    7  2  4 */ (n411 ? n337 : !n337);
assign n728  = /* LUT    5  2  1 */ (n5 ? (n11 ? 1'b1 : n9) : 1'b0);
assign n729  = /* LUT    5 14  3 */ n238;
assign n730  = /* LUT    4  6  4 */ n21;
assign n731  = /* LUT    7 14  5 */ (n18 ? (n15 ? n398 : n406) : n398);
assign n732  = /* LUT    6 10  1 */ (n174 ? (n170 ? (n300 ? !n46 : 1'b1) : (n300 ? n46 : 1'b0)) : (n170 ? (n300 ? n46 : 1'b0) : (n300 ? !n46 : 1'b1)));
assign n733  = /* LUT    8 10  3 */ n463;
assign n734  = /* LUT    6  2  6 */ (n334 ? (n333 ? (n335 ? 1'b0 : n84) : n335) : (n333 ? (n335 ? 1'b0 : !n84) : 1'b1));
assign n735  = /* LUT    9 11  1 */ (n47 ? n227 : n343);
assign n736  = /* LUT    5  3  2 */ (n163 ? (n56 ? (n243 ? 1'b1 : !n92) : (n243 ? !n92 : 1'b1)) : (n56 ? (n243 ? 1'b0 : n92) : (n243 ? n92 : 1'b0)));
assign n737  = /* LUT    7  3  4 */ (n418 ? (n413 ? 1'b1 : n242) : (n413 ? (n330 ? n242 : !n242) : n330));
assign n738  = /* LUT    5  6  7 */ (n271 ? (n94 ? n272 : 1'b0) : (n94 ? (n259 ? !n272 : n272) : !n259));
assign n739  = /* LUT    2  2  4 */ (n5 ? (n6 ? (n11 ? !n59 : n59) : 1'b0) : 1'b0);
assign n740  = /* LUT    7  6  6 */ (n68 ? (n149 ? (n169 ? 1'b0 : !n271) : (n169 ? 1'b1 : n271)) : (n169 ? !n271 : 1'b0));
assign n741  = /* LUT    8 13  4 */ n472;
assign n742  = /* LUT    8  5  0 */ (n442 ? (n13 ? 1'b1 : (n283 ? 1'b1 : n419)) : 1'b0);
assign n743  = /* LUT    6  5  7 */ (n352 ? (n354 ? (n351 ? n353 : !n353) : (n351 ? 1'b0 : n353)) : (n354 ? (n351 ? !n353 : 1'b0) : 1'b1));
assign n744  = /* LUT   11 11  7 */ n549;
assign n745  = /* LUT    5 10  1 */ (n307 ? (n78 ? n14 : 1'b1) : (n78 ? !n14 : 1'b0));
assign n746  = /* LUT    8  6  1 */ (n441 ? (n13 ? 1'b1 : (n283 ? 1'b1 : n419)) : 1'b0);
assign n747  = /* LUT    9 10  5 */ n512;
assign n748  = /* LUT    5 13  6 */ n229;
assign n749  = /* LUT    6  9  4 */ (n19 ? n297 : n287);
assign n750  = /* LUT    4  9  5 */ (n195 ? (n46 ? !n129 : 1'b1) : (n46 ? n129 : 1'b0));
assign n751  = /* LUT    8  9  6 */ n453;
assign n752  = /* LUT   11  7  0 */ n543;
assign n753  = /* LUT    2  6  6 */ n48;
assign n754  = /* LUT    5  2  5 */ (n152 ? (n241 ? !n246 : n246) : (n241 ? n246 : !n246));
assign n755  = /* LUT   11  8  1 */ (n14 ? !n419 : 1'b0);
assign n756  = /* LUT    1  8  0 */ !n19;
assign n757  = /* LUT    6 12  5 */ n314;
assign n758  = /* LUT    7  6  1 */ (n271 ? (n275 ? (n272 ? 1'b0 : !n68) : (n272 ? 1'b1 : n68)) : (n272 ? !n68 : 1'b0));
assign n759  = /* LUT    9  6  3 */ n495;
assign n760  = /* LUT    5  9  4 */ n213;
assign n761  = /* LUT    2  5  1 */ n65;
assign n762  = /* LUT    6  5  2 */ (n274 ? (n270 ? n267 : (n264 ? n267 : !n267)) : (n270 ? 1'b1 : n264));
assign n763  = /* LUT    4  5  3 */ (n17 ? (n174 ? n67 : !n67) : (n174 ? !n67 : n67));
assign n764  = /* LUT    8  5  4 */ (n435 ? 1'b0 : !n429);
assign n765  = /* LUT   11  3  7 */ (n537 ? 1'b0 : (n92 ? (n66 ? 1'b1 : n488) : 1'b1));
assign n766  = /* LUT    5 10  5 */ n211;
assign n767  = /* LUT    9 10  0 */ n506;
assign n768  = /* LUT    7 10  7 */ (n193 ? !n48 : n48);
assign n769  = /* LUT    5 13  1 */ n230;
assign n770  = /* LUT    7  2  3 */ (n329 ? (n344 ? (n415 ? 1'b0 : !n245) : (n415 ? 1'b1 : n245)) : (n344 ? (n415 ? 1'b1 : n245) : (n415 ? 1'b0 : !n245)));
assign n771  = /* LUT    4  9  0 */ (n19 ? n128 : n73);
assign n772  = /* LUT    8  9  1 */ (n452 ? (n18 ? (n15 ? !n461 : 1'b1) : 1'b1) : 1'b0);
assign n773  = /* LUT    4  6  3 */ n20;
assign n774  = /* LUT    9 13  1 */ n476;
assign n775  = /* LUT    5  5  2 */ (n149 ? (n265 ? !n16 : 1'b0) : (n265 ? (n16 ? !n258 : n258) : n258));
assign n776  = /* LUT    7  5  4 */ (n169 ? (n149 ? (n16 ? 1'b0 : !n184) : (n16 ? !n184 : 1'b0)) : (n149 ? (n16 ? 1'b0 : n184) : (n16 ? n184 : 1'b0)));
assign n777  = /* LUT    6 12  0 */ n317;
assign n778  = /* LUT    4 12  1 */ n145;
assign n779  = /* LUT    8  4  7 */ (n358 ? (n416 ? !n431 : n431) : (n416 ? n431 : !n431));
assign n780  = /* LUT    7  6  5 */ (n273 ? n359 : !n359);
assign n781  = /* LUT    7  9  1 */ n369;
assign n782  = /* LUT    8 13  3 */ n526;
assign n783  = /* LUT    9  9  3 */ n510;
assign n784  = /* LUT    6  5  6 */ (n352 ? (n351 ? (n354 ? 1'b0 : n353) : n354) : (n351 ? (n354 ? 1'b0 : !n353) : 1'b1));
assign n785  = /* LUT    4  5  7 */ (n116 ? (n25 ? n14 : 1'b1) : (n25 ? !n14 : 1'b0));
assign n786  = /* LUT   11  3  2 */ (n554 ? (n534 ? 1'b0 : !n538) : (n534 ? !n538 : 1'b0));
assign n787  = /* LUT    5 10  0 */ n206;
assign n788  = /* LUT    7 10  2 */ n377;
assign n789  = /* LUT    2  9  2 */ n77;
assign n790  = /* LUT    7  2  7 */ (n417 ? !n413 : 1'b0);
assign n791  = /* LUT    4  9  4 */ (n19 ? n129 : n126);
assign n792  = /* LUT    6  8  7 */ n308;
assign n793  = /* LUT    5  5  6 */ (n265 ? (n169 ? !n184 : n184) : 1'b0);
assign n794  = /* LUT    9  5  1 */ (n419 ? (n492 ? 1'b0 : (n66 ? !n185 : 1'b1)) : (n66 ? !n185 : 1'b1));
assign n795  = /* LUT    6 12  4 */ (n18 ? (n15 ? n320 : n319) : n320);
assign n796  = /* LUT    6  4  0 */ (n352 ? (n353 ? 1'b0 : !n351) : (n353 ? 1'b1 : n354));
assign n797  = /* LUT    8  4  2 */ (n426 ? 1'b0 : !n177);
assign n798  = /* LUT    7  6  0 */ (n384 ? (n149 ? (n278 ? !n286 : n286) : (n278 ? n286 : !n286)) : (n149 ? (n278 ? n286 : !n286) : (n278 ? !n286 : n286)));
assign n799  = /* LUT    2 13  4 */ n99;
assign n800  = /* LUT    5  9  3 */ (n195 ? !n78 : n78);
assign n801  = /* LUT    2  5  0 */ (n62 ? n63 : 1'b0);
assign n802  = /* LUT    7  9  5 */ n383;
assign n803  = /* LUT    4 13  6 */ n146;
assign n804  = /* LUT    4  5  2 */ n113;
assign n805  = /* LUT    8  5  3 */ (n433 ? (n13 ? 1'b1 : (n283 ? 1'b1 : n419)) : 1'b0);
assign n806  = /* LUT    9  9  7 */ (n504 ? (n530 ? (n250 ? 1'b1 : n14) : (n250 ? n14 : 1'b1)) : (n530 ? (n250 ? 1'b0 : !n14) : (n250 ? !n14 : 1'b0)));
assign n807  = /* LUT    6  5  1 */ (n274 ? (n270 ? (n264 ? !n267 : n267) : !n264) : (n270 ? 1'b0 : !n267));
assign n808  = /* LUT   11 11  1 */ n553;
assign n809  = /* LUT    5 12  4 */ (n223 ? (n96 ? (n214 ? !n39 : 1'b1) : (n214 ? 1'b1 : !n39)) : 1'b0);
assign n810  = /* LUT    7  1  6 */ (n326 ? 1'b0 : (n336 ? 1'b0 : (n334 ? n328 : 1'b1)));
assign n811  = /* LUT    7 12  6 */ n391;
assign n812  = /* LUT    4  8  3 */ (n194 ? (n46 ? !n127 : 1'b1) : (n46 ? n127 : 1'b0));
assign n813  = /* LUT   11  7  3 */ n290;
assign n814  = /* LUT   11 10  5 */ (n47 ? n499 : n425);
assign n815  = /* LUT    5  5  1 */ (n184 ? (n265 ? (n169 ? n266 : !n266) : n266) : (n265 ? n169 : 1'b0));
assign n816  = /* LUT    7 13  7 */ n388;
assign n817  = /* LUT    7  5  3 */ (n355 ? (n364 ? (n361 ? !n274 : 1'b0) : (n361 ? n274 : 1'b1)) : (n364 ? (n361 ? n274 : 1'b1) : (n361 ? !n274 : 1'b0)));
assign n818  = /* LUT    9  5  5 */ n491;
assign n819  = /* LUT    2  4  3 */ (n62 ? 1'b0 : (n57 ? 1'b0 : (n58 ? 1'b0 : !n63)));
assign n820  = /* LUT    6  4  4 */ (n5 ? !n156 : 1'b0);
assign n821  = /* LUT    8  4  6 */ (n358 ? (n422 ? !n431 : n431) : (n422 ? n431 : !n431));
assign n822  = /* LUT    6  7  6 */ n189;
assign n823  = /* LUT    4 13  1 */ n147;
assign n824  = /* LUT    7  9  0 */ (n19 ? !n371 : !n374);
assign n825  = /* LUT    9  6  6 */ n493;
assign n826  = /* LUT    9  9  2 */ n501;
assign n827  = /* LUT   11 11  5 */ (n552 ? (n345 ? n14 : 1'b1) : (n345 ? !n14 : 1'b0));
assign n830  = /* LUT    6 11  3 */ (n19 ? n312 : n289);
assign n831  = /* LUT    8 11  5 */ n467;
assign n832  = /* LUT    7  1  1 */ (n407 ? (n162 ? !n341 : n341) : 1'b0);
assign n833  = /* LUT    7 12  1 */ n390;
assign n834  = /* LUT    5  4  4 */ n165;
assign n835  = /* LUT    6  8  6 */ n376;
assign n836  = /* LUT    4  8  7 */ (n170 ? (n46 ? n74 : 1'b0) : (n46 ? !n74 : 1'b1));
assign n837  = /* LUT    7 13  2 */ n400;
assign n838  = /* LUT    9 13  4 */ n525;
assign n839  = /* LUT    5  5  5 */ (n173 ? (n168 ? (n262 ? !n123 : n123) : (n262 ? n123 : !n123)) : (n168 ? (n262 ? n123 : !n123) : (n262 ? !n123 : n123)));
assign n840  = /* LUT    2 12  2 */ n81;
assign n841  = /* LUT    7  5  7 */ (n362 ? (n356 ? n357 : !n357) : (n356 ? !n357 : n357));
assign n842  = /* LUT    8  4  1 */ (n428 ? (n437 ? 1'b0 : !n439) : (n437 ? !n438 : (n439 ? !n438 : n438)));
assign n843  = /* LUT    2  4  7 */ (n62 ? !n63 : n63);
assign n844  = /* LUT    6  7  1 */ (n18 ? (n15 ? 1'b1 : !n95) : (n15 ? !n191 : 1'b1));
assign n845  = /* LUT    8  7  3 */ (n367 ? (n13 ? 1'b0 : (n283 ? 1'b0 : !n419)) : 1'b0);
assign n846  = /* LUT    5  8  6 */ n203;
assign n847  = /* LUT    5 11  2 */ (n22 ? (n46 ? n216 : 1'b0) : (n46 ? !n216 : 1'b1));
assign n848  = /* LUT    4  4  5 */ n106;
assign n849  = /* LUT    8 11  0 */ n470;
assign n850  = /* LUT    6 11  7 */ (n19 ? n309 : n310);
assign n851  = /* LUT   11  9  3 */ n500;
assign n852  = /* LUT    5 12  3 */ (n228 ? (n18 ? (n15 ? !n51 : 1'b1) : 1'b1) : 1'b0);
assign n853  = /* LUT    2  8  0 */ (n19 ? n74 : n72);
assign n854  = /* LUT    6  8  1 */ (n284 ? (n18 ? (n15 ? !n319 : 1'b1) : 1'b1) : 1'b0);
assign n855  = /* LUT    7  1  5 */ (n335 ? (n84 ? (n334 ? 1'b0 : n333) : n334) : (n84 ? (n334 ? 1'b0 : !n333) : 1'b1));
assign n856  = /* LUT    4  8  2 */ (n193 ? (n194 ? (n77 ? n46 : 1'b0) : (n77 ? !n46 : 1'b1)) : (n194 ? (n77 ? !n46 : 1'b1) : (n77 ? n46 : 1'b0)));
assign n857  = /* LUT    7  4  1 */ n157;
assign n858  = /* LUT    8  8  3 */ n385;
assign n859  = /* LUT    7 12  5 */ n394;
assign n860  = /* LUT   11 10  4 */ (n47 ? n547 : n530);
assign n861  = /* LUT    5  5  0 */ (n182 ? (n263 ? (n122 ? n171 : !n171) : (n122 ? !n171 : n171)) : (n263 ? (n122 ? !n171 : n171) : (n122 ? n171 : !n171)));
assign n862  = /* LUT    7  5  2 */ (n93 ? (n356 ? n355 : !n355) : (n356 ? !n355 : n355));
assign n863  = /* LUT    4 11  3 */ (n39 ? n98 : (n24 ? n134 : !n134));
assign n864  = /* LUT    8 15  2 */ n485;
assign n865  = /* LUT    2  3  6 */ (n89 ? !n59 : n59);
assign n866  = /* LUT    6  7  5 */ n282;
assign n867  = /* LUT    8  7  7 */ n369;
assign n868  = /* LUT    4  4  0 */ n107;
assign n869  = /* LUT    5 11  6 */ (n22 ? (n46 ? n215 : 1'b0) : (n46 ? !n215 : 1'b1));
assign n870  = /* LUT    2  7  3 */ n28;
assign n871  = /* LUT    6 11  2 */ (n178 ? (n46 ? n312 : 1'b0) : (n46 ? !n312 : 1'b1));
assign n872  = /* LUT   11  6  2 */ (n528 ? (n13 ? 1'b0 : (n283 ? 1'b0 : !n419)) : 1'b0);
assign n873  = /* LUT    8 11  4 */ n221;
assign n874  = /* LUT   11  9  7 */ n387;
assign n875  = /* LUT    7  1  0 */ (n162 ? n341 : !n341);
assign n876  = /* LUT    7 12  0 */ n393;
assign n877  = /* LUT    5 12  7 */ n224;
assign n878  = /* LUT    9 12  2 */ n523;
assign n879  = /* LUT    4  8  6 */ (n170 ? (n195 ? (n31 ? !n46 : 1'b1) : (n31 ? n46 : 1'b0)) : (n195 ? (n31 ? n46 : 1'b0) : (n31 ? !n46 : 1'b1)));
assign n880  = /* LUT    6  3  3 */ (n249 ? (n239 ? n342 : 1'b1) : (n239 ? (n342 ? n247 : !n247) : !n247));
assign n881  = /* LUT    8  3  5 */ (n416 ? (n430 ? !n432 : n432) : (n430 ? n432 : !n432));
assign n882  = /* LUT    5  7  4 */ (n15 ? (n18 ? n191 : n199) : n191);
assign n885  = /* LUT    7  7  6 */ (n18 ? (n15 ? n95 : n199) : n95);
assign n886  = /* LUT    4 11  7 */ n139;
assign n887  = /* LUT    6  7  0 */ (n133 ? n291 : !n291);
assign n888  = /* LUT    8 15  6 */ n484;
assign n889  = /* LUT   11  5  5 */ n539;
assign n890  = /* LUT    7  8  7 */ (n39 ? n319 : (n378 ? n30 : !n30));
assign n891  = /* LUT    5 11  1 */ (n178 ? (n46 ? n219 : 1'b0) : (n46 ? !n219 : 1'b1));
assign n892  = /* LUT   11  6  6 */ n96;
assign n893  = /* LUT   11  9  2 */ n503;
assign n894  = /* LUT    7 12  4 */ (n39 ? n406 : (n385 ? n42 : !n42));
assign n895  = /* LUT    4  8  1 */ (n195 ? (n46 ? !n125 : 1'b1) : (n46 ? n125 : 1'b0));
assign n896  = /* LUT    7  4  0 */ (n425 ? (n260 ? (n346 ? 1'b1 : !n92) : (n346 ? !n92 : 1'b1)) : (n260 ? (n346 ? 1'b0 : n92) : (n346 ? n92 : 1'b0)));
assign n897  = /* LUT    8  3  0 */ (n447 ? (n430 ? !n432 : n432) : (n430 ? n432 : !n432));
assign n898  = /* LUT    8 14  0 */ n482;
assign n899  = /* LUT    6  3  7 */ (n109 ? (n256 ? (n348 ? n347 : !n347) : (n348 ? !n347 : n347)) : (n256 ? (n348 ? !n347 : n347) : (n348 ? n347 : !n347)));
assign n900  = /* LUT    6 14  7 */ n300;
assign n901  = /* LUT    6  6  3 */ (n279 ? (n169 ? n68 : !n68) : (n169 ? !n68 : n68));
assign n902  = /* LUT    9  4  7 */ (n488 ? (n527 ? !rst : 1'b0) : 1'b0);
assign n903  = /* LUT    7  7  1 */ n368;
assign n904  = /* LUT    9  7  3 */ n378;
assign n905  = /* LUT    2  3  5 */ (n88 ? !n10 : n10);
assign n906  = /* LUT    4  3  7 */ (n101 ? (n102 ? (n8 ? !n92 : 1'b1) : (n8 ? 1'b1 : !n92)) : (n102 ? (n8 ? n92 : 1'b0) : (n8 ? 1'b0 : n92)));
assign n907  = /* LUT    6  7  4 */ (n277 ? (n18 ? (n15 ? !n199 : 1'b1) : 1'b1) : 1'b0);
assign n908  = /* LUT    8  7  6 */ n29;
assign n909  = /* LUT   11 13  4 */ n100;
assign n910  = /* LUT   11  5  0 */ n542;
assign n911  = /* LUT    5  8  0 */ (n174 ? (n183 ? !n187 : n187) : (n183 ? n187 : !n187));
assign n912  = /* LUT    7  8  2 */ (n32 ? (n188 ? (n376 ? n46 : 1'b0) : (n376 ? !n46 : 1'b1)) : (n188 ? (n376 ? !n46 : 1'b1) : (n376 ? n46 : 1'b0)));
assign n913  = /* LUT    5 11  5 */ n210;
assign n914  = /* LUT    7 11  7 */ (n22 ? n345 : !n345);
assign n915  = /* LUT    4  7  4 */ n27;
assign n916  = /* LUT    6 10  5 */ (n19 ? n301 : n325);
assign n917  = /* LUT    6  2  1 */ (n335 ? (n334 ? (n84 ? n333 : !n333) : (n84 ? 1'b0 : n333)) : (n334 ? (n84 ? !n333 : 1'b0) : 1'b1));
assign n918  = /* LUT    6 13  1 */ n316;
assign n919  = /* LUT    8 10  7 */ n459;
assign n920  = /* LUT    8  2  3 */ (n421 ? (n414 ? (n413 ? 1'b0 : !n417) : (n413 ? 1'b1 : n417)) : (n413 ? !n417 : 1'b0));
assign n921  = /* LUT    9 11  5 */ n519;
assign n922  = /* LUT    5  3  6 */ (n92 ? (n158 ? (n167 ? !n8 : n8) : (n167 ? n8 : !n8)) : 1'b0);
assign n923  = /* LUT    2 10  3 */ n76;
assign n924  = /* LUT    5  6  2 */ (n272 ? (n94 ? (n271 ? n261 : !n261) : !n261) : (n94 ? n271 : 1'b1));
assign n925  = /* LUT    6  3  2 */ (n109 ? (n347 ? !n167 : n167) : (n347 ? n167 : !n167));
assign n926  = /* LUT    8  3  4 */ (n420 ? (n447 ? !n430 : n430) : (n447 ? n430 : !n430));
assign n927  = /* LUT    6  6  7 */ (n136 ? (n149 ? (n278 ? n286 : !n286) : (n278 ? !n286 : n286)) : (n149 ? (n278 ? !n286 : n286) : (n278 ? n286 : !n286)));
assign n928  = /* LUT   11 12  7 */ n234;
assign n929  = /* LUT   11  4  3 */ (n537 ? (n536 ? (n535 ? 1'b0 : !n534) : 1'b0) : 1'b0);
assign n930  = /* LUT    9  4  2 */ (n419 ? !n492 : 1'b0);
assign n931  = /* LUT    5  7  3 */ n281;
assign n935  = /* LUT    4 11  6 */ n140;
assign n936  = /* LUT    7  7  5 */ n366;
assign n937  = /* LUT    4  3  2 */ (n5 ? (n104 ? (n10 ? !n9 : 1'b0) : 1'b0) : 1'b0);
assign n938  = /* LUT    9  7  7 */ n496;
assign n939  = /* LUT    8  7  1 */ (n448 ? (n13 ? 1'b1 : (n283 ? 1'b1 : n419)) : 1'b0);
assign n940  = /* LUT    8  6  5 */ n378;
assign n941  = /* LUT    5 11  0 */ (n19 ? !n219 : !n217);
assign n942  = /* LUT    7 11  2 */ (n471 ? (n369 ? (n97 ? !n39 : 1'b1) : (n97 ? 1'b1 : !n39)) : 1'b0);
assign n943  = /* LUT    5 14  2 */ n236;
assign n944  = /* LUT    6 10  0 */ (n19 ? !n302 : !n306);
assign n945  = /* LUT   11  9  1 */ n546;
assign n946  = /* LUT    8 10  2 */ n462;
assign n947  = /* LUT    6  2  5 */ (n332 ? (n162 ? 1'b1 : n245) : (n162 ? 1'b0 : !n245));
assign n948  = /* LUT    8  2  7 */ (n257 ? (n91 ? (n416 ? n342 : !n342) : n416) : (n91 ? 1'b0 : n342));
assign n949  = /* LUT    9 11  0 */ (n47 ? n386 : n395);
assign n950  = /* LUT    5  3  1 */ (n9 ? (n11 ? (n10 ? 1'b1 : n59) : 1'b1) : (n11 ? 1'b1 : (n10 ? n59 : 1'b1)));
assign n951  = /* LUT    7  3  3 */ (n108 ? (n417 ? n242 : 1'b1) : (n330 ? (n417 ? 1'b1 : n242) : (n417 ? 1'b0 : !n242)));
assign n952  = /* LUT    4 10  0 */ (n18 ? 1'b0 : !n15);
assign n953  = /* LUT    9  3  5 */ (n2 ? (n66 ? 1'b1 : rst) : 1'b1);
assign n954  = /* LUT    2 10  7 */ n43;
assign n955  = /* LUT    5  6  6 */ (n23 ? (n171 ? (n179 ? n123 : !n123) : (n179 ? !n123 : n123)) : (n171 ? (n179 ? !n123 : n123) : (n179 ? n123 : !n123)));
assign n956  = /* LUT    6  3  6 */ (n91 ? (n239 ? n257 : 1'b1) : (n239 ? (n257 ? n247 : !n247) : !n247));
assign n957  = /* LUT    6  6  2 */ (n276 ? n273 : !n273);
assign n958  = /* LUT   11 12  2 */ n148;
assign n959  = /* LUT   11  4  7 */ (rst ? 1'b0 : (n115 ? 1'b1 : (n13 ? n434 : 1'b0)));
assign n960  = /* LUT    4 11  1 */ (n137 ? (n18 ? (n15 ? !n98 : 1'b1) : 1'b1) : 1'b0);
assign n961  = /* LUT    7  7  0 */ (n291 ? (n360 ? !n286 : n286) : (n360 ? n286 : !n286));
assign n962  = /* LUT    5  7  7 */ n190;
assign n963  = /* LUT    9  7  2 */ n529;
assign n964  = /* LUT    2  3  4 */ (n87 ? !n9 : n9);
assign n965  = /* LUT    2 14  4 */ n83;
assign n966  = /* LUT    4 14  6 */ (n18 ? (n15 ? n235 : n53) : n235);
assign n967  = /* LUT    8  6  0 */ (n449 ? (n13 ? 1'b1 : (n283 ? 1'b1 : n419)) : 1'b0);
assign n968  = /* LUT    6  9  3 */ (n200 ? (n46 ? n299 : 1'b0) : (n46 ? !n299 : 1'b1));
assign n969  = /* LUT    8  9  5 */ n456;
assign n970  = /* LUT    5  2  4 */ (n151 ? (n59 ? 1'b0 : (n10 ? !n11 : 1'b1)) : 1'b0);
assign n971  = /* LUT    5 14  6 */ n237;
assign n972  = /* LUT    4  6  7 */ n119;
assign n973  = /* LUT    6 10  4 */ (n15 ? (n18 ? n41 : n319) : n41);
assign n974  = /* LUT    6  2  0 */ (n257 ? (n239 ? !n91 : 1'b0) : (n239 ? (n91 ? n244 : !n244) : !n244));
assign n975  = /* LUT    8 10  6 */ n458;
assign n976  = /* LUT    8  2  2 */ (n409 ? (n340 ? (n418 ? 1'b1 : n108) : (n418 ? 1'b0 : !n108)) : (n340 ? (n418 ? 1'b0 : !n108) : (n418 ? 1'b1 : n108)));
assign n977  = /* LUT    9 11  4 */ n516;
assign n978  = /* LUT    5  3  5 */ (n5 ? !n10 : 1'b0);
assign n979  = /* LUT    7  3  7 */ (n92 ? (n167 ? (n155 ? n8 : !n8) : (n155 ? !n8 : n8)) : 1'b0);
assign n980  = /* LUT    5  6  1 */ (n275 ? (n94 ? !n68 : 1'b1) : (n94 ? (n68 ? !n261 : n261) : !n261));
assign n981  = /* LUT    4  2  0 */ (n9 ? !n10 : 1'b0);
assign n982  = /* LUT    8 13  7 */ n24;
assign n983  = /* LUT   11  4  2 */ (n537 ? (n536 ? (n535 ? n534 : 1'b0) : 1'b0) : 1'b0);
assign n984  = /* LUT    9  4  1 */ (n493 ? (n13 ? 1'b0 : (n283 ? 1'b0 : !n419)) : 1'b0);
assign n985  = /* LUT    1 12  5 */ !rst;
assign n986  = /* LUT    5  7  2 */ n176;
assign n987  = /* LUT    7  7  4 */ n367;
assign n988  = /* LUT    4  3  1 */ (n5 ? (n9 ? (n10 ? n104 : 1'b0) : 1'b0) : 1'b0);
assign n989  = /* LUT    4 14  1 */ n150;
assign n990  = /* LUT    9  7  6 */ n528;
assign n991  = /* LUT    5 10  4 */ n79;
assign n992  = /* LUT    5 13  0 */ (n18 ? (n15 ? 1'b1 : !n233) : (n15 ? !n231 : 1'b1));
assign n993  = /* LUT    8  6  4 */ (n69 ? (n13 ? 1'b0 : (n283 ? 1'b0 : !n419)) : 1'b0);
assign n994  = /* LUT    7  2  2 */ (n162 ? (n418 ? !n108 : 1'b1) : (n415 ? (n418 ? !n108 : 1'b1) : (n418 ? n108 : 1'b0)));
assign n995  = /* LUT    8  9  0 */ (n135 ? (n38 ? (n379 ? !n39 : 1'b1) : (n379 ? 1'b1 : !n39)) : 1'b0);
assign n996  = /* LUT    6  9  7 */ (n188 ? (n46 ? !n298 : 1'b1) : (n46 ? n298 : 1'b0));
assign n997  = /* LUT    4  6  2 */ n186;
assign n998  = /* LUT    8 10  1 */ (n18 ? (n15 ? n451 : n461) : n451);
assign n999  = /* LUT    6  2  4 */ (n84 ? (n333 ? (n335 ? 1'b1 : n334) : (n335 ? n334 : 1'b1)) : (n333 ? 1'b0 : n334));
assign n1000 = /* LUT    6 13  4 */ n323;
assign n1001 = /* LUT    8  2  6 */ (n414 ? n417 : !n417);
assign n1002 = /* LUT    5  3  0 */ (n10 ? (n11 ? (n9 ? 1'b0 : !n59) : 1'b0) : 1'b0);
assign n1003 = /* LUT    7  3  2 */ (rst ? 1'b1 : (n64 ? 1'b1 : n185));
assign n1004 = /* LUT    5  6  5 */ (n180 ? !n262 : n262);
assign n1005 = /* LUT    7  6  4 */ (n273 ? (n359 ? !n275 : n275) : (n359 ? n275 : !n275));
assign n1006 = /* LUT    8 13  2 */ n477;
assign n1007 = /* LUT    6  5  5 */ (n354 ? (n351 ? 1'b0 : !n353) : (n351 ? 1'b1 : n352));
assign n1008 = /* LUT   11  4  6 */ (n488 ? 1'b0 : (n13 ? 1'b0 : (n283 ? 1'b0 : !n5)));
assign n1009 = /* LUT    8  5  7 */ n221;
assign n1010 = /* LUT    9 10  3 */ n517;
assign n1011 = /* LUT    5 13  4 */ n225;
assign n1012 = /* LUT    6  9  2 */ (n19 ? n298 : n296);
assign n1013 = /* LUT    7  2  6 */ (n332 ? (n348 ? (n331 ? n341 : 1'b1) : (n331 ? !n341 : 1'b0)) : (n348 ? (n331 ? !n341 : 1'b0) : (n331 ? n341 : 1'b1)));
assign n1014 = /* LUT    4  9  3 */ (n195 ? (n46 ? !n128 : 1'b1) : (n46 ? n128 : 1'b0));
assign n1015 = /* LUT    8  9  4 */ n455;
assign n1016 = /* LUT   11  7  7 */ n544;
assign n1017 = /* LUT    5  2  3 */ (n10 ? 1'b0 : !n59);
assign n1018 = /* LUT    5 14  5 */ (n15 ? (n18 ? n218 : n53) : n218);
assign n1019 = /* LUT    7 14  7 */ n405;
assign n1020 = /* LUT    8  2  1 */ (n91 ? (n416 ? (n257 ? !n342 : n342) : !n342) : (n416 ? 1'b1 : !n257));
assign n1021 = /* LUT    6 12  3 */ n318;
assign n1022 = /* LUT    8 12  5 */ n469;
assign n1023 = /* LUT    5  6  0 */ (n168 ? (n180 ? (n262 ? !n123 : n123) : (n262 ? n123 : !n123)) : (n180 ? (n262 ? n123 : !n123) : (n262 ? !n123 : n123)));
assign n1024 = /* LUT    9  6  1 */ (rst ? 1'b0 : !n489);
assign n1025 = /* LUT    5  9  2 */ (n209 ? !n160 : n160);
assign n1026 = /* LUT    4 13  5 */ (n18 ? (n15 ? n233 : n51) : n233);
assign n1027 = /* LUT    8 13  6 */ (n15 ? (n18 ? n475 : n521) : n475);
assign n1028 = /* LUT    6  5  0 */ (n361 ? (n269 ? 1'b0 : !n267) : (n269 ? (n264 ? !n267 : n267) : !n264));
assign n1029 = /* LUT   11  4  1 */ (n487 ? (n115 ? 1'b0 : (n185 ? 1'b1 : !n66)) : 1'b0);
assign n1030 = /* LUT    7  9  4 */ n382;
assign n1031 = /* LUT    8  5  2 */ (n435 ? (n436 ? 1'b1 : n445) : (n436 ? n429 : (n445 ? n429 : !n429)));
assign n1032 = /* LUT    9  9  6 */ n509;
assign n1033 = /* LUT   11 11  0 */ n550;
assign n1034 = /* LUT    5 10  3 */ (n39 ? n53 : (n221 ? n293 : !n293));
assign n1035 = /* LUT    7 10  5 */ n40;
assign n1036 = /* LUT    8  6  3 */ (n440 ? (n13 ? 1'b1 : (n283 ? 1'b1 : n419)) : 1'b0);
assign n1037 = /* LUT    7  2  1 */ (n413 ? (n418 ? 1'b0 : (n417 ? n108 : !n108)) : (n418 ? (n417 ? n108 : !n108) : 1'b0));
assign n1038 = /* LUT    9 10  7 */ n508;
assign n1039 = /* LUT    2  9  5 */ n36;
assign n1040 = /* LUT    6  9  6 */ (n188 ? (n46 ? !n297 : 1'b1) : (n46 ? n297 : 1'b0));
assign n1041 = /* LUT    4  9  7 */ (n178 ? (n193 ? (n46 ? !n131 : 1'b1) : (n46 ? n131 : 1'b0)) : (n193 ? (n46 ? n131 : 1'b0) : (n46 ? !n131 : 1'b1)));
assign n1042 = /* LUT    4  6  1 */ n69;
assign n1043 = /* LUT    7 14  2 */ n404;
assign n1044 = /* LUT    5  2  7 */ (n241 ? (n246 ? (n153 ? n6 : 1'b1) : (n153 ? !n6 : 1'b0)) : (n246 ? (n153 ? !n6 : 1'b0) : (n153 ? n6 : 1'b1)));
assign n1045 = /* LUT    7 13  6 */ (n15 ? (n18 ? n402 : n406) : n402);
assign n1046 = /* LUT    8 12  0 */ (n473 ? (n18 ? (n15 ? !n521 : 1'b1) : 1'b1) : 1'b0);
assign n1047 = /* LUT    1  8  2 */ n31;
assign n1048 = /* LUT    6 12  7 */ n315;
assign n1049 = /* LUT    6  4  3 */ (n353 ? (n351 ? (n354 ? 1'b1 : n352) : (n354 ? n352 : 1'b1)) : (n351 ? 1'b0 : n352));
assign n1050 = /* LUT    8  4  5 */ (n428 ? 1'b0 : !n438);
assign n1051 = /* LUT    7  6  3 */ (n272 ? (n136 ? 1'b1 : !n271) : (n136 ? (n360 ? !n271 : n271) : !n360));
assign n1052 = /* LUT    8 13  1 */ (n18 ? (n15 ? 1'b1 : !n474) : (n15 ? !n475 : 1'b1));
assign n1053 = /* LUT    9  6  5 */ n494;
assign n1054 = /* LUT    5  9  6 */ n202;
assign n1055 = /* LUT    9  9  1 */ (n505 ? (n268 ? n14 : 1'b1) : (n268 ? !n14 : 1'b0));
assign n1056 = /* LUT    2  5  3 */ (n62 ? 1'b1 : (n57 ? (n63 ? 1'b1 : n58) : 1'b0));
assign n1057 = /* LUT    6  5  4 */ (n352 ? (n354 ? (n351 ? n353 : !n353) : n351) : (n354 ? n353 : (n351 ? n353 : !n353)));
assign n1058 = /* LUT    4  5  5 */ n110;
assign n1059 = /* LUT    8  5  6 */ (n444 ? (n427 ? 1'b0 : !n424) : (n427 ? !n446 : (n424 ? !n446 : n446)));
assign n1060 = /* LUT   11 11  4 */ n551;
assign n1064 = /* LUT    7 10  0 */ (n397 ? (n385 ? (n42 ? !n39 : 1'b1) : (n42 ? 1'b1 : !n39)) : 1'b0);
assign n1065 = /* LUT    5 10  7 */ n205;
assign n1066 = /* LUT    9 10  2 */ n511;
assign n1067 = /* LUT    7  2  5 */ (n408 ? n337 : !n337);
assign n1068 = /* LUT    4  9  2 */ (n178 ? (n187 ? (n36 ? n46 : 1'b0) : (n36 ? !n46 : 1'b1)) : (n187 ? (n36 ? !n46 : 1'b1) : (n36 ? n46 : 1'b0)));
assign n1069 = /* LUT    8  9  3 */ (n39 ? n461 : (n38 ? n379 : !n379));
assign n1070 = /* LUT    5  2  2 */ (n5 ? (n7 ? !n9 : n11) : 1'b0);
assign n1071 = /* LUT    7 13  1 */ (n396 ? (n18 ? (n15 ? !n406 : 1'b1) : 1'b1) : 1'b0);
assign n1072 = /* LUT    5  5  4 */ (n16 ? (n265 ? n149 : 1'b1) : (n265 ? (n149 ? n266 : !n266) : !n266));
assign n1073 = /* LUT    7  5  6 */ (n270 ? 1'b0 : !n269);
assign n1074 = /* LUT    6 12  2 */ n392;
assign n1075 = /* LUT    4 12  3 */ n144;
assign n1076 = /* LUT    8  4  0 */ (n422 ? (n437 ? 1'b1 : n439) : (n437 ? 1'b0 : !n439));
assign n1077 = /* LUT    2  4  6 */ !n62;
assign n1078 = /* LUT    6  4  7 */ (n354 ? (n353 ? (n352 ? 1'b0 : n351) : n352) : (n353 ? (n352 ? 1'b0 : !n351) : 1'b1));
assign n1079 = /* LUT    9  6  0 */ n490;
assign n1080 = /* LUT    5  9  1 */ (n178 ? n22 : !n22);
assign n1081 = /* LUT    7  6  7 */ n268;
assign n1082 = /* LUT    8 13  5 */ (n18 ? (n15 ? n474 : n521) : n474);
assign n1083 = /* LUT    7  9  3 */ n381;
assign n1084 = /* LUT    4  5  0 */ n112;
assign n1085 = /* LUT    8  5  1 */ (n490 ? (n13 ? 1'b0 : (n283 ? 1'b0 : !n419)) : 1'b0);
assign n1086 = /* LUT    9  9  5 */ n38;
assign n1087 = /* LUT   11  3  4 */ (n537 ? (n536 ? 1'b0 : !n538) : (n536 ? !n538 : 1'b0));
assign n1088 = /* LUT    7  2  0 */ (n411 ? (n408 ? (n337 ? 1'b0 : !n84) : 1'b0) : (n408 ? 1'b0 : (n337 ? !n84 : 1'b0)));
assign n1089 = /* LUT    7  1  4 */ (n335 ? (n334 ? (n84 ? n333 : !n333) : n84) : (n334 ? n333 : (n84 ? n333 : !n333)));
assign n1090 = /* LUT   11  7  1 */ n545;
assign n1091 = /* LUT    5  4  7 */ n164;
assign n1092 = /* LUT    7 13  5 */ n399;
assign n1093 = /* LUT    7  5  1 */ (n184 ? (n16 ? (n270 ? n269 : 1'b0) : (n270 ? !n269 : 1'b1)) : (n270 ? n269 : 1'b0));
assign n1094 = /* LUT    2 12  5 */ n80;
assign n1095 = /* LUT    6 12  6 */ n321;
assign n1096 = /* LUT    2  4  1 */ (rst ? 1'b1 : (n55 ? n61 : 1'b0));
assign n1097 = /* LUT    4 12  7 */ n143;
assign n1098 = /* LUT    6  4  2 */ (n353 ? (n354 ? !n351 : (n352 ? !n351 : 1'b1)) : (n354 ? 1'b0 : (n352 ? 1'b1 : !n351)));
assign n1099 = /* LUT    8  4  4 */ (n427 ? (n426 ? 1'b1 : n177) : (n426 ? n424 : (n177 ? n424 : !n424)));
assign n1100 = /* LUT   11  2  7 */ (n329 ? (n421 ? n331 : 1'b0) : (n421 ? !n331 : 1'b1));
assign n1101 = /* LUT    7  6  2 */ (n360 ? (n149 ? (n278 ? !n286 : n286) : (n278 ? n286 : !n286)) : (n149 ? (n278 ? n286 : !n286) : (n278 ? !n286 : n286)));
assign n1102 = /* LUT    9  6  4 */ n365;
assign n1103 = /* LUT    5  9  5 */ n37;
assign n1104 = /* LUT    9  9  0 */ n502;
assign n1105 = /* LUT    2  5  2 */ (n62 ? (n63 ? 1'b1 : n58) : (n63 ? n58 : 1'b1));
assign n1106 = /* LUT    7  9  7 */ n212;
assign n1107 = /* LUT    4  5  4 */ (n118 ? (n17 ? (n67 ? 1'b1 : n14) : (n67 ? n14 : 1'b1)) : (n17 ? (n67 ? 1'b0 : !n14) : (n67 ? !n14 : 1'b0)));
assign n1108 = /* LUT   11 11  3 */ n518;
assign n1109 = /* LUT    6 11  1 */ (n174 ? (n46 ? !n311 : 1'b1) : (n46 ? n311 : 1'b0));
assign n1110 = /* LUT    8 11  3 */ (n39 ? n521 : (n369 ? n97 : !n97));
assign n87   = /* CARRY  2  3  3 */ (1'b0 & n58) | ((1'b0 | n58) & n86);
assign n86   = /* CARRY  2  3  2 */ (1'b0 & n57) | ((1'b0 | n57) & n85);
assign n555  = /* CARRY 11  3  2 */ (1'b0 & n534) | ((1'b0 | n534) & n554);
assign n554  = /* CARRY 11  3  1 */ (1'b0 & n536) | ((1'b0 | n536) & n557);
assign n90   = /* CARRY  2  3  6 */ (1'b0 & n59) | ((1'b0 | n59) & n89);
assign n85   = /* CARRY  2  3  1 */ (1'b0 & n63) | ((1'b0 | n63) & n556);
assign n89   = /* CARRY  2  3  5 */ (1'b0 & n10) | ((1'b0 | n10) & n88);
assign n556  = /* CARRY  2  3  0 */ (n62 & 1'b0) | ((n62 | 1'b0) & n934);
assign n88   = /* CARRY  2  3  4 */ (1'b0 & n9) | ((1'b0 | n9) & n87);
assign n557  = /* CARRY 11  3  0 */ (n537 & 1'b0) | ((n537 | 1'b0) & n1063);
/* FF  5 12  6 */ always @(posedge clk) if (1'b1) n225 <= 1'b0 ? 1'b0 : n558;
/* FF  9 12  1 */ always @(posedge clk) if (1'b1) n234 <= 1'b0 ? 1'b0 : n559;
/* FF  2  8  3 */ always @(posedge clk) if (1'b1) n71 <= 1'b0 ? 1'b0 : n560;
/* FF  5  4  2 */ always @(posedge clk) if (1'b1) n163 <= 1'b0 ? 1'b0 : n561;
/* FF  6  8  4 */ always @(posedge clk) if (1'b1) n287 <= n4 ? 1'b1 : n562;
/* FF  4  8  5 */ always @(posedge clk) if (1'b1) n74 <= 1'b0 ? 1'b0 : n563;
/* FF  7 13  0 */ assign n396 = n564;
/* FF  5  5  3 */ assign n172 = n565;
/* FF  2 12  0 */ always @(posedge clk) if (1'b1) n80 <= 1'b0 ? 1'b0 : n566;
/* FF  7  5  5 */ assign n356 = n567;
/* FF  6 12  1 */ always @(posedge clk) if (1'b1) n315 <= 1'b0 ? 1'b0 : n568;
/* FF  4 12  2 */ always @(posedge clk) if (1'b1) n142 <= 1'b0 ? 1'b0 : n569;
/* FF  9  5  7 */ always @(posedge clk) if (1'b1) n491 <= 1'b0 ? 1'b0 : n570;
/* FF  8 15  5 */ always @(posedge clk) if (1'b1) n484 <= 1'b0 ? 1'b0 : n571;
/* FF  5  9  0 */ assign n136 = n572;
/* FF  7  9  2 */ always @(posedge clk) if (1'b1) n381 <= 1'b0 ? 1'b0 : n573;
/* FF  9  9  4 */ always @(posedge clk) if (1'b1) n505 <= 1'b0 ? 1'b0 : n574;
/* FF  5  8  4 */ assign n195 = n575;
/* FF  7  8  6 */ always @(posedge clk) if (1'b1) n376 <= 1'b0 ? 1'b0 : n576;
/* FF 11  3  3 */ always @(posedge clk) if (n486) n535 <= rst ? 1'b0 : n577;
/* FF  6 11  5 */ always @(posedge clk) if (1'b1) n312 <= 1'b0 ? 1'b0 : n578;
/* FF  8 11  7 */ always @(posedge clk) if (1'b1) n470 <= 1'b0 ? 1'b0 : n579;
/* FF  5 12  1 */ assign n192 = n580;
/* FF  7  1  3 */ assign n329 = n581;
/* FF  4  8  0 */ assign n30 = n582;
/* FF  9 12  5 */ always @(posedge clk) if (1'b1) n523 <= 1'b0 ? 1'b0 : n583;
/* FF  2  8  7 */ always @(posedge clk) if (1'b1) n72 <= 1'b0 ? 1'b0 : n584;
/* FF  5  4  6 */ always @(posedge clk) if (1'b1) n165 <= 1'b0 ? 1'b0 : n585;
/* FF  7 13  4 */ always @(posedge clk) if (1'b1) n399 <= 1'b0 ? 1'b0 : n586;
/* FF  7  5  0 */ assign n351 = n587;
/* FF  9 13  6 */ always @(posedge clk) if (1'b1) n525 <= 1'b0 ? 1'b0 : n588;
/* FF  5  5  7 */ always @(posedge clk) if (1'b1) n176 <= n2 ? 1'b0 : n589;
/* FF  4 12  6 */ always @(posedge clk) if (1'b1) n144 <= 1'b0 ? 1'b0 : n590;
/* FF  8  4  3 */ assign n421 = n591;
/* FF  8 15  0 */ always @(posedge clk) if (1'b1) n482 <= 1'b0 ? 1'b0 : n592;
/* FF  6  7  3 */ assign n279 = n593;
/* FF  8  7  5 */ assign n447 = n594;
/* FF  7  8  1 */ always @(posedge clk) if (1'b1) n372 <= 1'b0 ? 1'b0 : n595;
/* FF  9  8  3 */ always @(posedge clk) if (1'b1) n499 <= 1'b0 ? 1'b0 : n596;
/* FF  5 11  4 */ always @(posedge clk) if (1'b1) n217 <= 1'b0 ? 1'b0 : n597;
/* FF  4  4  7 */ always @(posedge clk) if (1'b1) n107 <= 1'b0 ? 1'b0 : n598;
/* FF  6 11  0 */ assign n97 = n599;
/* FF  8 11  2 */ always @(posedge clk) if (1'b1) n466 <= 1'b0 ? 1'b0 : n600;
/* FF  5 12  5 */ always @(posedge clk) if (1'b1) n224 <= 1'b0 ? 1'b0 : n601;
/* FF  6  8  3 */ assign n286 = n602;
/* FF  7  1  7 */ assign n333 = n603;
/* FF  4  8  4 */ always @(posedge clk) if (1'b1) n124 <= 1'b0 ? 1'b0 : n604;
/* FF  7 12  7 */ always @(posedge clk) if (1'b1) n394 <= 1'b0 ? 1'b0 : n605;
/* FF  6  3  1 */ assign n251 = n606;
/* FF  8  3  3 */ assign n162 = n607;
/* FF  1 10  5 */ always @(posedge clk) if (1'b1) n35 <= n2 ? 1'b1 : n608;
/* FF  6  6  6 */ assign n274 = n609;
/* FF  8  7  0 */ assign n443 = n610;
/* FF  6  7  7 */ always @(posedge clk) if (1'b1) n282 <= 1'b0 ? 1'b0 : n611;
/* FF  5  8  3 */ assign n194 = n612;
/* FF  7  8  5 */ always @(posedge clk) if (1'b1) n375 <= 1'b0 ? 1'b0 : n613;
/* FF  6 11  4 */ always @(posedge clk) if (1'b1) n311 <= 1'b0 ? 1'b0 : n614;
/* FF 11  6  4 */ assign n427 = n615;
/* FF 11  9  0 */ always @(posedge clk) if (1'b1) n546 <= 1'b0 ? 1'b0 : n616;
/* FF  5 12  0 */ assign n222 = n617;
/* FF  7  1  2 */ assign n328 = n618;
/* FF  7 12  2 */ always @(posedge clk) if (1'b1) n390 <= 1'b0 ? 1'b0 : n619;
/* FF  9 12  4 */ always @(posedge clk) if (1'b1) n522 <= 1'b0 ? 1'b0 : n620;
/* FF  2 11  2 */ always @(posedge clk) if (1'b1) n49 <= n4 ? 1'b0 : n621;
/* FF  6  3  5 */ assign n255 = n622;
/* FF  6  6  1 */ assign n270 = n623;
/* FF  8  3  7 */ assign n342 = n624;
/* FF  4 11  0 */ assign n137 = n625;
/* FF  9  4  5 */ always @(posedge clk) if (1'b1) n13 <= 1'b0 ? 1'b0 : n626;
/* FF  5  7  6 */ always @(posedge clk) if (1'b1) n116 <= 1'b0 ? 1'b0 : n627;
/* FF  9  7  1 */ always @(posedge clk) if (1'b1) n496 <= 1'b0 ? 1'b0 : n628;
/* FF  2  3  3 */ always @(posedge clk) if (1'b1) n58 <= n1 ? 1'b0 : n629;
/* FF  4  3  5 */ assign n104 = n630;
/* FF  6  7  2 */ assign n278 = n631;
/* FF  8  7  4 */ assign n446 = n632;
/* FF  7  8  0 */ always @(posedge clk) if (1'b1) n371 <= 1'b0 ? 1'b0 : n633;
/* FF  5  8  7 */ always @(posedge clk) if (1'b1) n197 <= 1'b0 ? 1'b0 : n634;
/* FF  5 11  3 */ always @(posedge clk) if (1'b1) n216 <= 1'b0 ? 1'b0 : n635;
/* FF  7 11  5 */ assign n48 = n636;
/* FF  8 11  1 */ always @(posedge clk) if (1'b1) n465 <= 1'b0 ? 1'b0 : n637;
/* FF  6 10  3 */ always @(posedge clk) if (1'b1) n303 <= 1'b0 ? 1'b0 : n638;
/* FF 11  9  4 */ always @(posedge clk) if (1'b1) n547 <= 1'b0 ? 1'b0 : n639;
/* FF  8 10  5 */ always @(posedge clk) if (1'b1) n461 <= 1'b0 ? 1'b0 : n640;
/* FF  9 11  3 */ always @(posedge clk) if (1'b1) n516 <= 1'b0 ? 1'b0 : n641;
/* FF  5  3  4 */ assign n67 = n642;
/* FF  2 10  1 */ always @(posedge clk) if (1'b1) n76 <= 1'b0 ? 1'b0 : n643;
/* FF  7  3  6 */ assign n12 = n644;
/* FF  4 10  3 */ assign n134 = n645;
/* FF  6  3  0 */ assign n250 = n646;
/* FF  8  3  2 */ assign n91 = n647;
/* FF  8 14  2 */ always @(posedge clk) if (1'b1) n480 <= 1'b0 ? 1'b0 : n648;
/* FF  6  6  5 */ assign n273 = n649;
/* FF  9  4  0 */ assign n487 = n650;
/* FF  5  7  1 */ assign n188 = n651;
/* FF  4 11  4 */ always @(posedge clk) if (1'b1) n140 <= 1'b0 ? 1'b0 : n652;
/* FF  7  7  3 */ always @(posedge clk) if (1'b1) n368 <= 1'b0 ? 1'b0 : n653;
/* FF  2  3  7 */ always @(posedge clk) if (1'b1) n11 <= n1 ? 1'b0 : n654;
/* FF 11  5  2 */ always @(posedge clk) if (1'b1) n240 <= 1'b0 ? 1'b0 : n655;
/* FF  5  8  2 */ assign n32 = n656;
/* FF  7  8  4 */ always @(posedge clk) if (1'b1) n374 <= 1'b0 ? 1'b0 : n657;
/* FF  9  8  6 */ always @(posedge clk) if (1'b1) n500 <= 1'b0 ? 1'b0 : n658;
/* FF  5 11  7 */ always @(posedge clk) if (1'b1) n220 <= 1'b0 ? 1'b0 : n659;
/* FF  4  7  6 */ always @(posedge clk) if (1'b1) n95 <= 1'b0 ? 1'b0 : n660;
/* FF  8 10  0 */ always @(posedge clk) if (1'b1) n458 <= 1'b0 ? 1'b0 : n661;
/* FF  6 10  7 */ always @(posedge clk) if (1'b1) n300 <= 1'b0 ? 1'b0 : n662;
/* FF  6  2  3 */ assign n244 = n663;
/* FF  8  2  5 */ assign n407 = n664;
/* FF  7  3  1 */ assign n346 = n665;
/* FF  9 11  7 */ always @(posedge clk) if (1'b1) n343 <= 1'b0 ? 1'b0 : n666;
/* FF  5  6  4 */ assign n182 = n667;
/* FF  4 10  7 */ assign n133 = n668;
/* FF  6  3  4 */ assign n254 = n669;
/* FF  6  6  0 */ assign n269 = n670;
/* FF  8  3  6 */ assign n418 = n671;
/* FF  8 14  6 */ always @(posedge clk) if (1'b1) n481 <= 1'b0 ? 1'b0 : n672;
/* FF 11  4  5 */ assign n92 = n673;
/* FF  9  4  4 */ always @(posedge clk) if (1'b1) n488 <= 1'b0 ? 1'b0 : n674;
/* FF  5  7  5 */ always @(posedge clk) if (1'b1) n186 <= 1'b0 ? 1'b0 : n675;
/* FF  9  7  0 */ always @(posedge clk) if (1'b1) n290 <= 1'b0 ? 1'b0 : n676;
/* FF  2 14  2 */ always @(posedge clk) if (1'b1) n83 <= 1'b0 ? 1'b0 : n677;
/* FF  7  7  7 */ always @(posedge clk) if (1'b1) n29 <= 1'b0 ? 1'b0 : n678;
/* FF  2  3  2 */ always @(posedge clk) if (1'b1) n57 <= n1 ? 1'b0 : n679;
/* FF  6  9  1 */ assign n293 = n680;
/* FF  8  6  7 */ always @(posedge clk) if (n5) n442 <= 1'b0 ? 1'b0 : n681;
/* FF  2  6  3 */ always @(posedge clk) if (1'b1) n21 <= n2 ? 1'b0 : n682;
/* FF  4  6  5 */ always @(posedge clk) if (1'b1) n46 <= 1'b0 ? 1'b0 : n683;
/* FF  6 10  2 */ always @(posedge clk) if (1'b1) n302 <= 1'b0 ? 1'b0 : n684;
/* FF  7 14  6 */ always @(posedge clk) if (1'b1) n405 <= 1'b0 ? 1'b0 : n685;
/* FF  8  2  0 */ assign n408 = n686;
/* FF  6  2  7 */ assign n248 = n687;
/* FF  6 13  7 */ always @(posedge clk) if (1'b1) n323 <= 1'b0 ? 1'b0 : n688;
/* FF 11  8  7 */ always @(posedge clk) if (1'b1) n545 <= n2 ? 1'b1 : n689;
/* FF  5  3  3 */ assign n158 = n690;
/* FF  7  3  5 */ assign n344 = n691;
/* FF  4 10  2 */ assign n42 = n692;
/* FF  8  3  1 */ assign n108 = n693;
/* FF  6  6  4 */ assign n272 = n694;
/* FF 11  4  0 */ assign n527 = n695;
/* FF  5  7  0 */ assign n187 = n696;
/* FF  7  7  2 */ always @(posedge clk) if (1'b1) n367 <= 1'b0 ? 1'b0 : n697;
/* FF  5 10  2 */ always @(posedge clk) if (1'b1) n207 <= 1'b0 ? 1'b0 : n698;
/* FF 11  5  1 */ always @(posedge clk) if (1'b1) n66 <= 1'b0 ? 1'b0 : n699;
/* FF  8  6  2 */ assign n438 = n700;
/* FF  9 10  6 */ always @(posedge clk) if (1'b1) n512 <= 1'b0 ? 1'b0 : n701;
/* FF  5 13  7 */ always @(posedge clk) if (1'b1) n233 <= 1'b0 ? 1'b0 : n702;
/* FF  6  9  5 */ always @(posedge clk) if (1'b1) n297 <= 1'b0 ? 1'b0 : n703;
/* FF  4  9  6 */ always @(posedge clk) if (1'b1) n132 <= 1'b0 ? 1'b0 : n704;
/* FF  8  9  7 */ always @(posedge clk) if (1'b1) n457 <= 1'b0 ? 1'b0 : n705;
/* FF  6  1  1 */ assign n239 = n706;
/* FF  4  6  0 */ always @(posedge clk) if (1'b1) \d_out[7]  <= 1'b0 ? 1'b0 : n707;
/* FF  5  2  6 */ assign n154 = n708;
/* FF  6 10  6 */ always @(posedge clk) if (1'b1) n306 <= 1'b0 ? 1'b0 : n709;
/* FF  6  2  2 */ assign n243 = n710;
/* FF  8  2  4 */ assign n411 = n711;
/* FF 11  8  2 */ always @(posedge clk) if (1'b1) n544 <= n2 ? 1'b1 : n712;
/* FF  7  3  0 */ assign n345 = n713;
/* FF  9 11  6 */ always @(posedge clk) if (1'b1) n519 <= 1'b0 ? 1'b0 : n714;
/* FF  5  3  7 */ always @(posedge clk) if (1'b1) \d_out[5]  <= 1'b0 ? 1'b0 : n715;
/* FF  5  6  3 */ assign n181 = n716;
/* FF  2  2  0 */ assign n55 = n717;
/* FF  6  5  3 */ assign n263 = n718;
/* FF 11  4  4 */ assign n434 = n719;
/* FF  8  5  5 */ assign n431 = n720;
/* FF  5 10  6 */ always @(posedge clk) if (1'b1) n210 <= 1'b0 ? 1'b0 : n721;
/* FF  5 13  2 */ always @(posedge clk) if (1'b1) n230 <= 1'b0 ? 1'b0 : n722;
/* FF  6  9  0 */ assign n284 = n723;
/* FF  8  6  6 */ always @(posedge clk) if (n5) n441 <= 1'b0 ? 1'b0 : n724;
/* FF  4  9  1 */ always @(posedge clk) if (1'b1) n127 <= 1'b0 ? 1'b0 : n725;
/* FF  8  9  2 */ assign n452 = n726;
/* FF  7  2  4 */ assign n334 = n727;
/* FF  5  2  1 */ assign n151 = n728;
/* FF  5 14  3 */ always @(posedge clk) if (1'b1) n236 <= 1'b0 ? 1'b0 : n729;
/* FF  4  6  4 */ always @(posedge clk) if (1'b1) n120 <= 1'b0 ? 1'b0 : n730;
/* FF  7 14  5 */ always @(posedge clk) if (1'b1) n404 <= 1'b0 ? 1'b0 : n731;
/* FF  6 10  1 */ always @(posedge clk) if (1'b1) n301 <= 1'b0 ? 1'b0 : n732;
/* FF  8 10  3 */ always @(posedge clk) if (1'b1) n460 <= 1'b0 ? 1'b0 : n733;
/* FF  6  2  6 */ assign n247 = n734;
/* FF  9 11  1 */ assign \d_out[0]  = n735;
/* FF  5  3  2 */ assign n157 = n736;
/* FF  7  3  4 */ assign n348 = n737;
/* FF  5  6  7 */ assign n23 = n738;
/* FF  2  2  4 */ assign n56 = n739;
/* FF  7  6  6 */ assign n364 = n740;
/* FF  8 13  4 */ always @(posedge clk) if (1'b1) n475 <= 1'b0 ? 1'b0 : n741;
/* FF  8  5  0 */ assign n428 = n742;
/* FF  6  5  7 */ assign n267 = n743;
/* FF 11 11  7 */ always @(posedge clk) if (1'b1) n552 <= 1'b0 ? 1'b0 : n744;
/* FF  5 10  1 */ always @(posedge clk) if (1'b1) n206 <= 1'b0 ? 1'b0 : n745;
/* FF  8  6  1 */ assign n437 = n746;
/* FF  9 10  5 */ always @(posedge clk) if (1'b1) n511 <= 1'b0 ? 1'b0 : n747;
/* FF  5 13  6 */ always @(posedge clk) if (1'b1) n232 <= 1'b0 ? 1'b0 : n748;
/* FF  6  9  4 */ always @(posedge clk) if (1'b1) n296 <= 1'b0 ? 1'b0 : n749;
/* FF  4  9  5 */ always @(posedge clk) if (1'b1) n131 <= 1'b0 ? 1'b0 : n750;
/* FF  8  9  6 */ always @(posedge clk) if (1'b1) n456 <= 1'b0 ? 1'b0 : n751;
/* FF 11  7  0 */ always @(posedge clk) if (1'b1) n528 <= 1'b0 ? 1'b0 : n752;
/* FF  2  6  6 */ always @(posedge clk) if (1'b1) n20 <= n2 ? 1'b1 : n753;
/* FF  5  2  5 */ assign n105 = n754;
/* FF 11  8  1 */ assign n2 = n755;
/* FF  1  8  0 */ assign n4 = n756;
/* FF  6 12  5 */ always @(posedge clk) if (1'b1) n319 <= 1'b0 ? 1'b0 : n757;
/* FF  7  6  1 */ assign n362 = n758;
/* FF  9  6  3 */ always @(posedge clk) if (1'b1) n38 <= 1'b0 ? 1'b0 : n759;
/* FF  5  9  4 */ always @(posedge clk) if (1'b1) n202 <= 1'b0 ? 1'b0 : n760;
/* FF  2  5  1 */ always @(posedge clk) if (1'b1) n19 <= n66 ? 1'b0 : n761;
/* FF  6  5  2 */ assign n122 = n762;
/* FF  4  5  3 */ always @(posedge clk) if (1'b1) \d_out[6]  <= 1'b0 ? 1'b0 : n763;
/* FF  8  5  4 */ assign n430 = n764;
/* FF 11  3  7 */ always @(posedge clk) if (n486) n537 <= rst ? 1'b0 : n765;
/* FF  5 10  5 */ always @(posedge clk) if (1'b1) n209 <= 1'b0 ? 1'b0 : n766;
/* FF  9 10  0 */ always @(posedge clk) if (1'b1) n508 <= 1'b0 ? 1'b0 : n767;
/* FF  7 10  7 */ always @(posedge clk) if (1'b1) n386 <= 1'b0 ? 1'b0 : n768;
/* FF  5 13  1 */ always @(posedge clk) if (1'b1) n229 <= 1'b0 ? 1'b0 : n769;
/* FF  7  2  3 */ assign n339 = n770;
/* FF  4  9  0 */ always @(posedge clk) if (1'b1) n126 <= 1'b0 ? 1'b0 : n771;
/* FF  8  9  1 */ assign n135 = n772;
/* FF  4  6  3 */ always @(posedge clk) if (1'b1) n119 <= 1'b0 ? 1'b0 : n773;
/* FF  9 13  1 */ always @(posedge clk) if (1'b1) n524 <= 1'b0 ? 1'b0 : n774;
/* FF  5  5  2 */ assign n171 = n775;
/* FF  7  5  4 */ assign n355 = n776;
/* FF  6 12  0 */ always @(posedge clk) if (1'b1) n314 <= 1'b0 ? 1'b0 : n777;
/* FF  4 12  1 */ always @(posedge clk) if (1'b1) n98 <= 1'b0 ? 1'b0 : n778;
/* FF  8  4  7 */ assign n413 = n779;
/* FF  7  6  5 */ assign n184 = n780;
/* FF  7  9  1 */ always @(posedge clk) if (1'b1) n380 <= 1'b0 ? 1'b0 : n781;
/* FF  8 13  3 */ always @(posedge clk) if (1'b1) n474 <= 1'b0 ? 1'b0 : n782;
/* FF  9  9  3 */ always @(posedge clk) if (1'b1) n504 <= 1'b0 ? 1'b0 : n783;
/* FF  6  5  6 */ assign n266 = n784;
/* FF  4  5  7 */ always @(posedge clk) if (1'b1) n114 <= 1'b0 ? 1'b0 : n785;
/* FF 11  3  2 */ always @(posedge clk) if (n486) n534 <= rst ? 1'b0 : n786;
/* FF  5 10  0 */ always @(posedge clk) if (1'b1) n205 <= 1'b0 ? 1'b0 : n787;
/* FF  7 10  2 */ always @(posedge clk) if (1'b1) n79 <= 1'b0 ? 1'b0 : n788;
/* FF  2  9  2 */ always @(posedge clk) if (1'b1) n70 <= n4 ? 1'b1 : n789;
/* FF  7  2  7 */ assign n340 = n790;
/* FF  4  9  4 */ always @(posedge clk) if (1'b1) n130 <= 1'b0 ? 1'b0 : n791;
/* FF  6  8  7 */ always @(posedge clk) if (1'b1) n289 <= n4 ? 1'b0 : n792;
/* FF  5  5  6 */ assign n175 = n793;
/* FF  9  5  1 */ assign n489 = n794;
/* FF  6 12  4 */ always @(posedge clk) if (1'b1) n318 <= 1'b0 ? 1'b0 : n795;
/* FF  6  4  0 */ assign n94 = n796;
/* FF  8  4  2 */ assign n416 = n797;
/* FF  7  6  0 */ assign n169 = n798;
/* FF  2 13  4 */ always @(posedge clk) if (1'b1) n51 <= 1'b0 ? 1'b0 : n799;
/* FF  5  9  3 */ always @(posedge clk) if (1'b1) \d_out[4]  <= 1'b0 ? 1'b0 : n800;
/* FF  2  5  0 */ assign n65 = n801;
/* FF  7  9  5 */ always @(posedge clk) if (1'b1) n37 <= 1'b0 ? 1'b0 : n802;
/* FF  4 13  6 */ always @(posedge clk) if (1'b1) n147 <= 1'b0 ? 1'b0 : n803;
/* FF  4  5  2 */ always @(posedge clk) if (1'b1) n17 <= 1'b0 ? 1'b0 : n804;
/* FF  8  5  3 */ assign n426 = n805;
/* FF  9  9  7 */ always @(posedge clk) if (1'b1) n387 <= 1'b0 ? 1'b0 : n806;
/* FF  6  5  1 */ assign n262 = n807;
/* FF 11 11  1 */ always @(posedge clk) if (1'b1) n549 <= 1'b0 ? 1'b0 : n808;
/* FF  5 12  4 */ assign n149 = n809;
/* FF  7  1  6 */ assign n332 = n810;
/* FF  7 12  6 */ always @(posedge clk) if (1'b1) n393 <= 1'b0 ? 1'b0 : n811;
/* FF  4  8  3 */ always @(posedge clk) if (1'b1) n77 <= 1'b0 ? 1'b0 : n812;
/* FF 11  7  3 */ always @(posedge clk) if (1'b1) n542 <= 1'b0 ? 1'b0 : n813;
/* FF 11 10  5 */ assign \d_out[2]  = n814;
/* FF  5  5  1 */ assign n168 = n815;
/* FF  7 13  7 */ always @(posedge clk) if (1'b1) n402 <= 1'b0 ? 1'b0 : n816;
/* FF  7  5  3 */ assign n353 = n817;
/* FF  9  5  5 */ always @(posedge clk) if (1'b1) n490 <= 1'b0 ? 1'b0 : n818;
/* FF  2  4  3 */ assign n61 = n819;
/* FF  6  4  4 */ assign n260 = n820;
/* FF  8  4  6 */ assign n257 = n821;
/* FF  6  7  6 */ always @(posedge clk) if (1'b1) n198 <= 1'b0 ? 1'b0 : n822;
/* FF  4 13  1 */ always @(posedge clk) if (1'b1) n99 <= 1'b0 ? 1'b0 : n823;
/* FF  7  9  0 */ assign n379 = n824;
/* FF  9  6  6 */ always @(posedge clk) if (1'b1) n221 <= 1'b0 ? 1'b0 : n825;
/* FF  9  9  2 */ always @(posedge clk) if (1'b1) n503 <= 1'b0 ? 1'b0 : n826;
/* FF 11 11  5 */ always @(posedge clk) if (1'b1) n551 <= 1'b0 ? 1'b0 : n827;
/* FF 11  3  1 */ assign n828 = n829;
/* FF  6 11  3 */ always @(posedge clk) if (1'b1) n310 <= 1'b0 ? 1'b0 : n830;
/* FF  8 11  5 */ always @(posedge clk) if (1'b1) n469 <= 1'b0 ? 1'b0 : n831;
/* FF  7  1  1 */ assign n327 = n832;
/* FF  7 12  1 */ always @(posedge clk) if (1'b1) n389 <= 1'b0 ? 1'b0 : n833;
/* FF  5  4  4 */ always @(posedge clk) if (1'b1) n164 <= 1'b0 ? 1'b0 : n834;
/* FF  6  8  6 */ always @(posedge clk) if (1'b1) n288 <= n4 ? 1'b0 : n835;
/* FF  4  8  7 */ always @(posedge clk) if (1'b1) n125 <= 1'b0 ? 1'b0 : n836;
/* FF  7 13  2 */ always @(posedge clk) if (1'b1) n398 <= 1'b0 ? 1'b0 : n837;
/* FF  9 13  4 */ always @(posedge clk) if (1'b1) n521 <= 1'b0 ? 1'b0 : n838;
/* FF  5  5  5 */ assign n174 = n839;
/* FF  2 12  2 */ always @(posedge clk) if (1'b1) n50 <= 1'b0 ? 1'b0 : n840;
/* FF  7  5  7 */ assign n354 = n841;
/* FF  8  4  1 */ assign n358 = n842;
/* FF  2  4  7 */ always @(posedge clk) if (1'b1) n63 <= n1 ? 1'b0 : n843;
/* FF  6  7  1 */ assign n277 = n844;
/* FF  8  7  3 */ assign n445 = n845;
/* FF  5  8  6 */ always @(posedge clk) if (1'b1) n196 <= 1'b0 ? 1'b0 : n846;
/* FF  5 11  2 */ always @(posedge clk) if (1'b1) n215 <= 1'b0 ? 1'b0 : n847;
/* FF  4  4  5 */ always @(posedge clk) if (1'b1) n101 <= 1'b0 ? 1'b0 : n848;
/* FF  8 11  0 */ always @(posedge clk) if (1'b1) n464 <= 1'b0 ? 1'b0 : n849;
/* FF  6 11  7 */ always @(posedge clk) if (1'b1) n313 <= 1'b0 ? 1'b0 : n850;
/* FF 11  9  3 */ always @(posedge clk) if (1'b1) n212 <= 1'b0 ? 1'b0 : n851;
/* FF  5 12  3 */ assign n223 = n852;
/* FF  2  8  0 */ always @(posedge clk) if (1'b1) n34 <= 1'b0 ? 1'b0 : n853;
/* FF  6  8  1 */ assign n285 = n854;
/* FF  7  1  5 */ assign n331 = n855;
/* FF  4  8  2 */ always @(posedge clk) if (1'b1) n33 <= 1'b0 ? 1'b0 : n856;
/* FF  7  4  1 */ always @(posedge clk) if (1'b1) n350 <= n2 ? 1'b0 : n857;
/* FF  8  8  3 */ always @(posedge clk) if (n5) n450 <= 1'b0 ? 1'b0 : n858;
/* FF  7 12  5 */ always @(posedge clk) if (1'b1) n392 <= 1'b0 ? 1'b0 : n859;
/* FF 11 10  4 */ assign \d_out[1]  = n860;
/* FF  5  5  0 */ assign n170 = n861;
/* FF  7  5  2 */ assign n352 = n862;
/* FF  4 11  3 */ always @(posedge clk) if (1'b1) n139 <= 1'b0 ? 1'b0 : n863;
/* FF  8 15  2 */ always @(posedge clk) if (1'b1) n483 <= 1'b0 ? 1'b0 : n864;
/* FF  2  3  6 */ always @(posedge clk) if (1'b1) n59 <= n1 ? 1'b0 : n865;
/* FF  6  7  5 */ always @(posedge clk) if (1'b1) n281 <= 1'b0 ? 1'b0 : n866;
/* FF  8  7  7 */ always @(posedge clk) if (n5) n449 <= 1'b0 ? 1'b0 : n867;
/* FF  4  4  0 */ always @(posedge clk) if (1'b1) n106 <= 1'b0 ? 1'b0 : n868;
/* FF  5 11  6 */ always @(posedge clk) if (1'b1) n219 <= 1'b0 ? 1'b0 : n869;
/* FF  2  7  3 */ always @(posedge clk) if (1'b1) n27 <= 1'b0 ? 1'b0 : n870;
/* FF  6 11  2 */ always @(posedge clk) if (1'b1) n309 <= 1'b0 ? 1'b0 : n871;
/* FF 11  6  2 */ assign n424 = n872;
/* FF  8 11  4 */ always @(posedge clk) if (1'b1) n468 <= 1'b0 ? 1'b0 : n873;
/* FF 11  9  7 */ always @(posedge clk) if (1'b1) n548 <= 1'b0 ? 1'b0 : n874;
/* FF  7  1  0 */ assign n326 = n875;
/* FF  7 12  0 */ always @(posedge clk) if (1'b1) n388 <= 1'b0 ? 1'b0 : n876;
/* FF  5 12  7 */ always @(posedge clk) if (1'b1) n226 <= 1'b0 ? 1'b0 : n877;
/* FF  9 12  2 */ always @(posedge clk) if (1'b1) n148 <= 1'b0 ? 1'b0 : n878;
/* FF  4  8  6 */ always @(posedge clk) if (1'b1) n75 <= 1'b0 ? 1'b0 : n879;
/* FF  6  3  3 */ assign n253 = n880;
/* FF  8  3  5 */ assign n249 = n881;
/* FF  5  7  4 */ always @(posedge clk) if (1'b1) n28 <= 1'b0 ? 1'b0 : n882;
/* FF  2  3  1 */ assign n883 = n884;
/* FF  7  7  6 */ always @(posedge clk) if (1'b1) n370 <= 1'b0 ? 1'b0 : n885;
/* FF  4 11  7 */ always @(posedge clk) if (1'b1) n141 <= 1'b0 ? 1'b0 : n886;
/* FF  6  7  0 */ assign n276 = n887;
/* FF  8 15  6 */ always @(posedge clk) if (1'b1) n485 <= 1'b0 ? 1'b0 : n888;
/* FF 11  5  5 */ always @(posedge clk) if (1'b1) n540 <= 1'b0 ? 1'b0 : n889;
/* FF  7  8  7 */ always @(posedge clk) if (1'b1) n377 <= 1'b0 ? 1'b0 : n890;
/* FF  5 11  1 */ always @(posedge clk) if (1'b1) n45 <= 1'b0 ? 1'b0 : n891;
/* FF 11  6  6 */ always @(posedge clk) if (n5) n541 <= 1'b0 ? 1'b0 : n892;
/* FF 11  9  2 */ always @(posedge clk) if (1'b1) n425 <= 1'b0 ? 1'b0 : n893;
/* FF  7 12  4 */ always @(posedge clk) if (1'b1) n391 <= 1'b0 ? 1'b0 : n894;
/* FF  4  8  1 */ always @(posedge clk) if (1'b1) n31 <= 1'b0 ? 1'b0 : n895;
/* FF  7  4  0 */ assign n268 = n896;
/* FF  8  3  0 */ assign n415 = n897;
/* FF  8 14  0 */ always @(posedge clk) if (1'b1) n479 <= 1'b0 ? 1'b0 : n898;
/* FF  6  3  7 */ assign n8 = n899;
/* FF  6 14  7 */ always @(posedge clk) if (1'b1) n325 <= n4 ? 1'b0 : n900;
/* FF  6  6  3 */ assign n16 = n901;
/* FF  9  4  7 */ always @(posedge clk) if (1'b1) n283 <= 1'b0 ? 1'b0 : n902;
/* FF  7  7  1 */ always @(posedge clk) if (1'b1) n366 <= 1'b0 ? 1'b0 : n903;
/* FF  9  7  3 */ always @(posedge clk) if (1'b1) n497 <= 1'b0 ? 1'b0 : n904;
/* FF  2  3  5 */ always @(posedge clk) if (1'b1) n10 <= n1 ? 1'b0 : n905;
/* FF  4  3  7 */ assign n25 = n906;
/* FF  6  7  4 */ assign n280 = n907;
/* FF  8  7  6 */ always @(posedge clk) if (n5) n448 <= 1'b0 ? 1'b0 : n908;
/* FF 11 13  4 */ always @(posedge clk) if (1'b1) n526 <= 1'b0 ? 1'b0 : n909;
/* FF 11  5  0 */ always @(posedge clk) if (1'b1) n539 <= 1'b0 ? 1'b0 : n910;
/* FF  5  8  0 */ assign n193 = n911;
/* FF  7  8  2 */ always @(posedge clk) if (1'b1) n373 <= 1'b0 ? 1'b0 : n912;
/* FF  5 11  5 */ always @(posedge clk) if (1'b1) n218 <= 1'b0 ? 1'b0 : n913;
/* FF  7 11  7 */ always @(posedge clk) if (1'b1) n227 <= 1'b0 ? 1'b0 : n914;
/* FF  4  7  4 */ always @(posedge clk) if (1'b1) n121 <= 1'b0 ? 1'b0 : n915;
/* FF  6 10  5 */ always @(posedge clk) if (1'b1) n305 <= 1'b0 ? 1'b0 : n916;
/* FF  6  2  1 */ assign n242 = n917;
/* FF  6 13  1 */ always @(posedge clk) if (1'b1) n322 <= 1'b0 ? 1'b0 : n918;
/* FF  8 10  7 */ always @(posedge clk) if (1'b1) n463 <= 1'b0 ? 1'b0 : n919;
/* FF  8  2  3 */ assign n410 = n920;
/* FF  9 11  5 */ always @(posedge clk) if (1'b1) n518 <= 1'b0 ? 1'b0 : n921;
/* FF  5  3  6 */ assign n160 = n922;
/* FF  2 10  3 */ always @(posedge clk) if (1'b1) n40 <= 1'b0 ? 1'b0 : n923;
/* FF  5  6  2 */ assign n180 = n924;
/* FF  6  3  2 */ assign n252 = n925;
/* FF  8  3  4 */ assign n417 = n926;
/* FF  6  6  7 */ assign n275 = n927;
/* FF 11 12  7 */ always @(posedge clk) if (1'b1) n553 <= 1'b0 ? 1'b0 : n928;
/* FF 11  4  3 */ assign n492 = n929;
/* FF  9  4  2 */ assign n115 = n930;
/* FF  5  7  3 */ always @(posedge clk) if (1'b1) n190 <= 1'b0 ? 1'b0 : n931;
/* FF  2  3  0 */ assign n932 = n933;
/* FF  4 11  6 */ always @(posedge clk) if (1'b1) n82 <= 1'b0 ? 1'b0 : n935;
/* FF  7  7  5 */ always @(posedge clk) if (1'b1) n199 <= 1'b0 ? 1'b0 : n936;
/* FF  4  3  2 */ assign n103 = n937;
/* FF  9  7  7 */ always @(posedge clk) if (1'b1) n498 <= 1'b0 ? 1'b0 : n938;
/* FF  8  7  1 */ assign n444 = n939;
/* FF  8  6  5 */ always @(posedge clk) if (n5) n440 <= 1'b0 ? 1'b0 : n940;
/* FF  5 11  0 */ assign n214 = n941;
/* FF  7 11  2 */ assign n360 = n942;
/* FF  5 14  2 */ always @(posedge clk) if (1'b1) n235 <= 1'b0 ? 1'b0 : n943;
/* FF  6 10  0 */ assign n292 = n944;
/* FF 11  9  1 */ always @(posedge clk) if (1'b1) n530 <= 1'b0 ? 1'b0 : n945;
/* FF  8 10  2 */ always @(posedge clk) if (1'b1) n451 <= 1'b0 ? 1'b0 : n946;
/* FF  6  2  5 */ assign n246 = n947;
/* FF  8  2  7 */ assign n412 = n948;
/* FF  9 11  0 */ assign \d_out[3]  = n949;
/* FF  5  3  1 */ assign n156 = n950;
/* FF  7  3  3 */ assign n347 = n951;
/* FF  4 10  0 */ assign n39 = n952;
/* FF  9  3  5 */ assign n486 = n953;
/* FF  2 10  7 */ always @(posedge clk) if (1'b1) n41 <= 1'b0 ? 1'b0 : n954;
/* FF  5  6  6 */ assign n22 = n955;
/* FF  6  3  6 */ assign n256 = n956;
/* FF  6  6  2 */ assign n271 = n957;
/* FF 11 12  2 */ always @(posedge clk) if (1'b1) n324 <= 1'b0 ? 1'b0 : n958;
/* FF 11  4  7 */ always @(posedge clk) if (1'b1) n419 <= 1'b0 ? 1'b0 : n959;
/* FF  4 11  1 */ assign n138 = n960;
/* FF  7  7  0 */ assign n359 = n961;
/* FF  5  7  7 */ always @(posedge clk) if (1'b1) n191 <= 1'b0 ? 1'b0 : n962;
/* FF  9  7  2 */ always @(posedge clk) if (1'b1) n493 <= 1'b0 ? 1'b0 : n963;
/* FF  2  3  4 */ always @(posedge clk) if (1'b1) n9 <= n1 ? 1'b0 : n964;
/* FF  2 14  4 */ always @(posedge clk) if (1'b1) n53 <= 1'b0 ? 1'b0 : n965;
/* FF  4 14  6 */ always @(posedge clk) if (1'b1) n150 <= 1'b0 ? 1'b0 : n966;
/* FF  8  6  0 */ assign n436 = n967;
/* FF  6  9  3 */ always @(posedge clk) if (1'b1) n295 <= 1'b0 ? 1'b0 : n968;
/* FF  8  9  5 */ always @(posedge clk) if (1'b1) n455 <= 1'b0 ? 1'b0 : n969;
/* FF  5  2  4 */ assign n153 = n970;
/* FF  5 14  6 */ always @(posedge clk) if (1'b1) n238 <= 1'b0 ? 1'b0 : n971;
/* FF  4  6  7 */ always @(posedge clk) if (1'b1) n69 <= 1'b0 ? 1'b0 : n972;
/* FF  6 10  4 */ always @(posedge clk) if (1'b1) n304 <= 1'b0 ? 1'b0 : n973;
/* FF  6  2  0 */ assign n241 = n974;
/* FF  8 10  6 */ always @(posedge clk) if (1'b1) n462 <= 1'b0 ? 1'b0 : n975;
/* FF  8  2  2 */ assign n84 = n976;
/* FF  9 11  4 */ always @(posedge clk) if (1'b1) n517 <= 1'b0 ? 1'b0 : n977;
/* FF  5  3  5 */ assign n159 = n978;
/* FF  7  3  7 */ assign n349 = n979;
/* FF  5  6  1 */ assign n179 = n980;
/* FF  4  2  0 */ assign n6 = n981;
/* FF  8 13  7 */ always @(posedge clk) if (1'b1) n478 <= 1'b0 ? 1'b0 : n982;
/* FF 11  4  2 */ assign n185 = n983;
/* FF  9  4  1 */ assign n177 = n984;
/* FF  1 12  5 */ always @(posedge clk) if (n60) d_vld <= 1'b0 ? 1'b0 : n985;
/* FF  5  7  2 */ always @(posedge clk) if (1'b1) n189 <= 1'b0 ? 1'b0 : n986;
/* FF  7  7  4 */ always @(posedge clk) if (1'b1) n369 <= 1'b0 ? 1'b0 : n987;
/* FF  4  3  1 */ assign n102 = n988;
/* FF  4 14  1 */ always @(posedge clk) if (1'b1) n54 <= 1'b0 ? 1'b0 : n989;
/* FF  9  7  6 */ always @(posedge clk) if (1'b1) n96 <= 1'b0 ? 1'b0 : n990;
/* FF  5 10  4 */ always @(posedge clk) if (1'b1) n43 <= 1'b0 ? 1'b0 : n991;
/* FF  5 13  0 */ assign n228 = n992;
/* FF  8  6  4 */ assign n439 = n993;
/* FF  7  2  2 */ assign n338 = n994;
/* FF  8  9  0 */ assign n291 = n995;
/* FF  6  9  7 */ always @(posedge clk) if (1'b1) n299 <= 1'b0 ? 1'b0 : n996;
/* FF  4  6  2 */ always @(posedge clk) if (1'b1) n118 <= 1'b0 ? 1'b0 : n997;
/* FF  8 10  1 */ always @(posedge clk) if (1'b1) n459 <= 1'b0 ? 1'b0 : n998;
/* FF  6  2  4 */ assign n245 = n999;
/* FF  6 13  4 */ always @(posedge clk) if (1'b1) n307 <= 1'b0 ? 1'b0 : n1000;
/* FF  8  2  6 */ assign n341 = n1001;
/* FF  5  3  0 */ assign n64 = n1002;
/* FF  7  3  2 */ assign n1 = n1003;
/* FF  5  6  5 */ assign n183 = n1004;
/* FF  7  6  4 */ assign n361 = n1005;
/* FF  8 13  2 */ always @(posedge clk) if (1'b1) n100 <= 1'b0 ? 1'b0 : n1006;
/* FF  6  5  5 */ assign n265 = n1007;
/* FF 11  4  6 */ assign n14 = n1008;
/* FF  8  5  7 */ always @(posedge clk) if (n5) n433 <= 1'b0 ? 1'b0 : n1009;
/* FF  9 10  3 */ always @(posedge clk) if (1'b1) n510 <= 1'b0 ? 1'b0 : n1010;
/* FF  5 13  4 */ always @(posedge clk) if (1'b1) n231 <= 1'b0 ? 1'b0 : n1011;
/* FF  6  9  2 */ always @(posedge clk) if (1'b1) n294 <= 1'b0 ? 1'b0 : n1012;
/* FF  7  2  6 */ assign n167 = n1013;
/* FF  4  9  3 */ always @(posedge clk) if (1'b1) n129 <= 1'b0 ? 1'b0 : n1014;
/* FF  8  9  4 */ always @(posedge clk) if (1'b1) n454 <= 1'b0 ? 1'b0 : n1015;
/* FF 11  7  7 */ always @(posedge clk) if (1'b1) n543 <= 1'b0 ? 1'b0 : n1016;
/* FF  5  2  3 */ assign n7 = n1017;
/* FF  5 14  5 */ always @(posedge clk) if (1'b1) n237 <= 1'b0 ? 1'b0 : n1018;
/* FF  7 14  7 */ always @(posedge clk) if (1'b1) n406 <= 1'b0 ? 1'b0 : n1019;
/* FF  8  2  1 */ assign n409 = n1020;
/* FF  6 12  3 */ always @(posedge clk) if (1'b1) n317 <= 1'b0 ? 1'b0 : n1021;
/* FF  8 12  5 */ always @(posedge clk) if (1'b1) n472 <= 1'b0 ? 1'b0 : n1022;
/* FF  5  6  0 */ assign n178 = n1023;
/* FF  9  6  1 */ always @(posedge clk) if (1'b1) n5 <= 1'b0 ? 1'b0 : n1024;
/* FF  5  9  2 */ assign n78 = n1025;
/* FF  4 13  5 */ always @(posedge clk) if (1'b1) n146 <= 1'b0 ? 1'b0 : n1026;
/* FF  8 13  6 */ always @(posedge clk) if (1'b1) n477 <= 1'b0 ? 1'b0 : n1027;
/* FF  6  5  0 */ assign n123 = n1028;
/* FF 11  4  1 */ assign n538 = n1029;
/* FF  7  9  4 */ always @(posedge clk) if (1'b1) n213 <= 1'b0 ? 1'b0 : n1030;
/* FF  8  5  2 */ assign n420 = n1031;
/* FF  9  9  6 */ always @(posedge clk) if (1'b1) n507 <= 1'b0 ? 1'b0 : n1032;
/* FF 11 11  0 */ always @(posedge clk) if (1'b1) n532 <= 1'b0 ? 1'b0 : n1033;
/* FF  5 10  3 */ always @(posedge clk) if (1'b1) n208 <= 1'b0 ? 1'b0 : n1034;
/* FF  7 10  5 */ always @(posedge clk) if (1'b1) n385 <= 1'b0 ? 1'b0 : n1035;
/* FF  8  6  3 */ assign n435 = n1036;
/* FF  7  2  1 */ assign n337 = n1037;
/* FF  9 10  7 */ always @(posedge clk) if (1'b1) n513 <= 1'b0 ? 1'b0 : n1038;
/* FF  2  9  5 */ always @(posedge clk) if (1'b1) n73 <= n4 ? 1'b1 : n1039;
/* FF  6  9  6 */ always @(posedge clk) if (1'b1) n298 <= 1'b0 ? 1'b0 : n1040;
/* FF  4  9  7 */ always @(posedge clk) if (1'b1) n36 <= 1'b0 ? 1'b0 : n1041;
/* FF  4  6  1 */ always @(posedge clk) if (1'b1) n24 <= 1'b0 ? 1'b0 : n1042;
/* FF  7 14  2 */ always @(posedge clk) if (1'b1) n403 <= 1'b0 ? 1'b0 : n1043;
/* FF  5  2  7 */ assign n155 = n1044;
/* FF  7 13  6 */ always @(posedge clk) if (1'b1) n401 <= 1'b0 ? 1'b0 : n1045;
/* FF  8 12  0 */ assign n471 = n1046;
/* FF  1  8  2 */ always @(posedge clk) if (1'b1) n26 <= n4 ? 1'b0 : n1047;
/* FF  6 12  7 */ always @(posedge clk) if (1'b1) n321 <= 1'b0 ? 1'b0 : n1048;
/* FF  6  4  3 */ assign n259 = n1049;
/* FF  8  4  5 */ assign n423 = n1050;
/* FF  7  6  3 */ assign n363 = n1051;
/* FF  8 13  1 */ assign n473 = n1052;
/* FF  9  6  5 */ always @(posedge clk) if (1'b1) n495 <= 1'b0 ? 1'b0 : n1053;
/* FF  5  9  6 */ always @(posedge clk) if (1'b1) n204 <= 1'b0 ? 1'b0 : n1054;
/* FF  9  9  1 */ always @(posedge clk) if (1'b1) n502 <= 1'b0 ? 1'b0 : n1055;
/* FF  2  5  3 */ always @(posedge clk) if (1'b1) n15 <= n66 ? 1'b1 : n1056;
/* FF  6  5  4 */ assign n264 = n1057;
/* FF  4  5  5 */ always @(posedge clk) if (1'b1) n113 <= 1'b0 ? 1'b0 : n1058;
/* FF  8  5  6 */ assign n432 = n1059;
/* FF 11 11  4 */ always @(posedge clk) if (1'b1) n550 <= 1'b0 ? 1'b0 : n1060;
/* FF 11  3  0 */ assign n1061 = n1062;
/* FF  7 10  0 */ assign n384 = n1064;
/* FF  5 10  7 */ always @(posedge clk) if (1'b1) n211 <= 1'b0 ? 1'b0 : n1065;
/* FF  9 10  2 */ always @(posedge clk) if (1'b1) n509 <= 1'b0 ? 1'b0 : n1066;
/* FF  7  2  5 */ assign n335 = n1067;
/* FF  4  9  2 */ always @(posedge clk) if (1'b1) n128 <= 1'b0 ? 1'b0 : n1068;
/* FF  8  9  3 */ always @(posedge clk) if (1'b1) n453 <= 1'b0 ? 1'b0 : n1069;
/* FF  5  2  2 */ assign n152 = n1070;
/* FF  7 13  1 */ assign n397 = n1071;
/* FF  5  5  4 */ assign n173 = n1072;
/* FF  7  5  6 */ assign n357 = n1073;
/* FF  6 12  2 */ always @(posedge clk) if (1'b1) n316 <= 1'b0 ? 1'b0 : n1074;
/* FF  4 12  3 */ always @(posedge clk) if (1'b1) n143 <= 1'b0 ? 1'b0 : n1075;
/* FF  8  4  0 */ assign n414 = n1076;
/* FF  2  4  6 */ always @(posedge clk) if (1'b1) n62 <= n1 ? 1'b0 : n1077;
/* FF  6  4  7 */ assign n261 = n1078;
/* FF  9  6  0 */ always @(posedge clk) if (1'b1) n378 <= 1'b0 ? 1'b0 : n1079;
/* FF  5  9  1 */ assign n200 = n1080;
/* FF  7  6  7 */ always @(posedge clk) if (1'b1) n365 <= n2 ? 1'b1 : n1081;
/* FF  8 13  5 */ always @(posedge clk) if (1'b1) n476 <= 1'b0 ? 1'b0 : n1082;
/* FF  7  9  3 */ always @(posedge clk) if (1'b1) n382 <= 1'b0 ? 1'b0 : n1083;
/* FF  4  5  0 */ always @(posedge clk) if (1'b1) n110 <= 1'b0 ? 1'b0 : n1084;
/* FF  8  5  1 */ assign n429 = n1085;
/* FF  9  9  5 */ always @(posedge clk) if (1'b1) n506 <= 1'b0 ? 1'b0 : n1086;
/* FF 11  3  4 */ always @(posedge clk) if (n486) n536 <= rst ? 1'b0 : n1087;
/* FF  7  2  0 */ assign n336 = n1088;
/* FF  7  1  4 */ assign n330 = n1089;
/* FF 11  7  1 */ always @(posedge clk) if (1'b1) n529 <= 1'b0 ? 1'b0 : n1090;
/* FF  5  4  7 */ always @(posedge clk) if (1'b1) n166 <= 1'b0 ? 1'b0 : n1091;
/* FF  7 13  5 */ always @(posedge clk) if (1'b1) n400 <= 1'b0 ? 1'b0 : n1092;
/* FF  7  5  1 */ assign n93 = n1093;
/* FF  2 12  5 */ always @(posedge clk) if (1'b1) n81 <= 1'b0 ? 1'b0 : n1094;
/* FF  6 12  6 */ always @(posedge clk) if (1'b1) n320 <= 1'b0 ? 1'b0 : n1095;
/* FF  2  4  1 */ assign n60 = n1096;
/* FF  4 12  7 */ always @(posedge clk) if (1'b1) n145 <= 1'b0 ? 1'b0 : n1097;
/* FF  6  4  2 */ assign n258 = n1098;
/* FF  8  4  4 */ assign n422 = n1099;
/* FF 11  2  7 */ assign n109 = n1100;
/* FF  7  6  2 */ assign n68 = n1101;
/* FF  9  6  4 */ always @(posedge clk) if (1'b1) n494 <= 1'b0 ? 1'b0 : n1102;
/* FF  5  9  5 */ always @(posedge clk) if (1'b1) n203 <= 1'b0 ? 1'b0 : n1103;
/* FF  9  9  0 */ always @(posedge clk) if (1'b1) n501 <= 1'b0 ? 1'b0 : n1104;
/* FF  2  5  2 */ always @(posedge clk) if (1'b1) n18 <= n66 ? 1'b1 : n1105;
/* FF  7  9  7 */ always @(posedge clk) if (1'b1) n383 <= 1'b0 ? 1'b0 : n1106;
/* FF  4  5  4 */ always @(posedge clk) if (1'b1) n112 <= 1'b0 ? 1'b0 : n1107;
/* FF 11 11  3 */ always @(posedge clk) if (1'b1) n395 <= 1'b0 ? 1'b0 : n1108;
/* FF  6 11  1 */ always @(posedge clk) if (1'b1) n308 <= 1'b0 ? 1'b0 : n1109;
/* FF  8 11  3 */ always @(posedge clk) if (1'b1) n467 <= 1'b0 ? 1'b0 : n1110;

endmodule

