// Reading file './modified_aes_blif/Modified_aes.asc'..

module chip (input clk, input rst, input select, output d_vld, output \d_out[5] , output \d_out[7] , output \d_out[6] , output \d_out[4] , output \d_out[1] , output \d_out[0] , output \d_out[2] , output \d_out[3] );

wire n1;
// (0, 0, 'glb_netwk_0')
// (1, 7, 'lutff_global/s_r')
// (2, 3, 'glb2local_2')
// (2, 3, 'local_g0_6')
// (2, 3, 'lutff_3/in_3')
// (4, 6, 'lutff_global/s_r')
// (5, 1, 'neigh_op_tnr_2')
// (5, 2, 'neigh_op_rgt_2')
// (5, 3, 'neigh_op_bnr_2')
// (5, 7, 'lutff_global/s_r')
// (6, 1, 'neigh_op_top_2')
// (6, 1, 'sp4_r_v_b_16')
// (6, 2, 'lutff_2/out')
// (6, 2, 'sp4_r_v_b_5')
// (6, 3, 'neigh_op_bot_2')
// (7, 0, 'fabout')
// (7, 0, 'local_g1_0')
// (7, 0, 'span4_vert_16')
// (7, 1, 'neigh_op_tnl_2')
// (7, 1, 'sp4_v_b_16')
// (7, 2, 'neigh_op_lft_2')
// (7, 2, 'sp4_v_b_5')
// (7, 3, 'neigh_op_bnl_2')
// (9, 6, 'lutff_global/s_r')
// (11, 4, 'lutff_global/s_r')
// (11, 10, 'lutff_global/s_r')

wire clk;
// (0, 0, 'glb_netwk_3')
// (0, 5, 'span4_vert_t_14')
// (0, 6, 'span4_vert_b_14')
// (0, 7, 'span4_vert_b_10')
// (0, 8, 'io_1/D_IN_0')
// (0, 8, 'io_1/PAD')
// (0, 8, 'span4_vert_b_6')
// (0, 9, 'fabout')
// (0, 9, 'local_g1_2')
// (0, 9, 'span4_vert_b_2')
// (1, 3, 'lutff_global/clk')
// (1, 5, 'lutff_global/clk')
// (1, 6, 'lutff_global/clk')
// (1, 7, 'lutff_global/clk')
// (1, 7, 'neigh_op_tnl_2')
// (1, 7, 'neigh_op_tnl_6')
// (1, 8, 'neigh_op_lft_2')
// (1, 8, 'neigh_op_lft_6')
// (1, 9, 'neigh_op_bnl_2')
// (1, 9, 'neigh_op_bnl_6')
// (2, 2, 'lutff_global/clk')
// (2, 3, 'lutff_global/clk')
// (2, 5, 'lutff_global/clk')
// (2, 6, 'lutff_global/clk')
// (2, 7, 'lutff_global/clk')
// (2, 8, 'lutff_global/clk')
// (2, 9, 'lutff_global/clk')
// (2, 10, 'lutff_global/clk')
// (2, 11, 'lutff_global/clk')
// (2, 14, 'lutff_global/clk')
// (4, 2, 'lutff_global/clk')
// (4, 3, 'lutff_global/clk')
// (4, 4, 'lutff_global/clk')
// (4, 5, 'lutff_global/clk')
// (4, 6, 'lutff_global/clk')
// (4, 7, 'lutff_global/clk')
// (4, 8, 'lutff_global/clk')
// (4, 9, 'lutff_global/clk')
// (4, 10, 'lutff_global/clk')
// (4, 11, 'lutff_global/clk')
// (4, 12, 'lutff_global/clk')
// (4, 14, 'lutff_global/clk')
// (5, 4, 'lutff_global/clk')
// (5, 5, 'lutff_global/clk')
// (5, 6, 'lutff_global/clk')
// (5, 7, 'lutff_global/clk')
// (5, 8, 'lutff_global/clk')
// (5, 9, 'lutff_global/clk')
// (5, 10, 'lutff_global/clk')
// (5, 11, 'lutff_global/clk')
// (5, 12, 'lutff_global/clk')
// (5, 13, 'lutff_global/clk')
// (5, 14, 'lutff_global/clk')
// (6, 3, 'lutff_global/clk')
// (6, 6, 'lutff_global/clk')
// (6, 9, 'lutff_global/clk')
// (6, 10, 'lutff_global/clk')
// (6, 11, 'lutff_global/clk')
// (6, 12, 'lutff_global/clk')
// (6, 13, 'lutff_global/clk')
// (7, 6, 'lutff_global/clk')
// (7, 9, 'lutff_global/clk')
// (7, 10, 'lutff_global/clk')
// (7, 11, 'lutff_global/clk')
// (7, 12, 'lutff_global/clk')
// (7, 13, 'lutff_global/clk')
// (7, 14, 'lutff_global/clk')
// (7, 15, 'lutff_global/clk')
// (8, 9, 'lutff_global/clk')
// (8, 10, 'lutff_global/clk')
// (8, 11, 'lutff_global/clk')
// (8, 12, 'lutff_global/clk')
// (8, 13, 'lutff_global/clk')
// (8, 14, 'lutff_global/clk')
// (9, 3, 'lutff_global/clk')
// (9, 4, 'lutff_global/clk')
// (9, 5, 'lutff_global/clk')
// (9, 6, 'lutff_global/clk')
// (9, 7, 'lutff_global/clk')
// (9, 8, 'lutff_global/clk')
// (9, 9, 'lutff_global/clk')
// (9, 10, 'lutff_global/clk')
// (9, 11, 'lutff_global/clk')
// (9, 12, 'lutff_global/clk')
// (9, 13, 'lutff_global/clk')
// (9, 14, 'lutff_global/clk')
// (11, 3, 'lutff_global/clk')
// (11, 4, 'lutff_global/clk')
// (11, 5, 'lutff_global/clk')
// (11, 6, 'lutff_global/clk')
// (11, 7, 'lutff_global/clk')
// (11, 8, 'lutff_global/clk')
// (11, 9, 'lutff_global/clk')
// (11, 10, 'lutff_global/clk')
// (11, 11, 'lutff_global/clk')
// (11, 12, 'lutff_global/clk')
// (11, 13, 'lutff_global/clk')
// (12, 9, 'lutff_global/clk')
// (12, 10, 'lutff_global/clk')
// (12, 11, 'lutff_global/clk')
// (12, 12, 'lutff_global/clk')

wire n3;
// (0, 0, 'glb_netwk_4')
// (5, 13, 'neigh_op_tnr_6')
// (5, 14, 'neigh_op_rgt_6')
// (5, 14, 'sp4_r_v_b_44')
// (5, 15, 'neigh_op_bnr_6')
// (5, 15, 'sp4_r_v_b_33')
// (5, 16, 'sp4_r_v_b_20')
// (6, 13, 'neigh_op_top_6')
// (6, 13, 'sp4_v_t_44')
// (6, 14, 'lutff_6/out')
// (6, 14, 'sp4_v_b_44')
// (6, 15, 'neigh_op_bot_6')
// (6, 15, 'sp4_v_b_33')
// (6, 16, 'sp4_v_b_20')
// (6, 17, 'fabout')
// (6, 17, 'local_g0_1')
// (6, 17, 'span4_vert_9')
// (7, 13, 'neigh_op_tnl_6')
// (7, 14, 'neigh_op_lft_6')
// (7, 15, 'neigh_op_bnl_6')
// (8, 14, 'lutff_global/s_r')
// (9, 7, 'lutff_global/s_r')
// (9, 10, 'lutff_global/s_r')
// (11, 11, 'lutff_global/s_r')
// (12, 9, 'lutff_global/s_r')
// (12, 12, 'lutff_global/s_r')

reg n4 = 0;
// (0, 0, 'glb_netwk_5')
// (3, 1, 'neigh_op_tnr_7')
// (3, 1, 'sp4_r_v_b_43')
// (3, 2, 'neigh_op_rgt_7')
// (3, 2, 'sp4_r_v_b_30')
// (3, 3, 'neigh_op_bnr_7')
// (3, 3, 'sp4_r_v_b_19')
// (3, 4, 'sp4_r_v_b_6')
// (4, 0, 'span4_horz_r_3')
// (4, 0, 'span4_vert_43')
// (4, 1, 'neigh_op_top_7')
// (4, 1, 'sp4_v_b_43')
// (4, 2, 'lutff_7/out')
// (4, 2, 'sp4_v_b_30')
// (4, 3, 'glb2local_0')
// (4, 3, 'glb2local_3')
// (4, 3, 'local_g0_4')
// (4, 3, 'local_g0_7')
// (4, 3, 'lutff_0/in_0')
// (4, 3, 'lutff_5/in_2')
// (4, 3, 'neigh_op_bot_7')
// (4, 3, 'sp4_v_b_19')
// (4, 4, 'sp4_v_b_6')
// (4, 6, 'glb2local_1')
// (4, 6, 'local_g0_5')
// (4, 6, 'lutff_0/in_3')
// (4, 6, 'lutff_4/in_3')
// (5, 0, 'span4_horz_r_7')
// (5, 1, 'neigh_op_tnl_7')
// (5, 2, 'neigh_op_lft_7')
// (5, 3, 'neigh_op_bnl_7')
// (5, 4, 'lutff_global/cen')
// (5, 5, 'lutff_global/cen')
// (6, 0, 'fabout')
// (6, 0, 'local_g0_3')
// (6, 0, 'span4_horz_r_11')
// (6, 3, 'lutff_global/cen')
// (6, 6, 'lutff_global/cen')
// (7, 0, 'span4_horz_r_15')
// (7, 5, 'glb2local_0')
// (7, 5, 'glb2local_1')
// (7, 5, 'local_g0_4')
// (7, 5, 'local_g0_5')
// (7, 5, 'lutff_2/in_3')
// (7, 5, 'lutff_4/in_3')
// (7, 5, 'lutff_7/in_3')
// (7, 6, 'glb2local_1')
// (7, 6, 'local_g0_5')
// (7, 6, 'lutff_2/in_3')
// (7, 6, 'lutff_6/in_3')
// (7, 6, 'lutff_global/cen')
// (8, 0, 'span4_horz_l_15')

wire n5;
// (0, 0, 'glb_netwk_6')
// (0, 6, 'span4_horz_31')
// (0, 6, 'span4_vert_t_13')
// (0, 7, 'span4_vert_b_13')
// (0, 8, 'fabout')
// (0, 8, 'local_g0_1')
// (0, 8, 'span4_vert_b_9')
// (0, 9, 'span4_vert_b_5')
// (0, 10, 'span4_vert_b_1')
// (1, 5, 'lutff_global/s_r')
// (1, 5, 'neigh_op_tnr_2')
// (1, 6, 'neigh_op_rgt_2')
// (1, 6, 'sp4_h_r_42')
// (1, 7, 'neigh_op_bnr_2')
// (2, 5, 'lutff_global/s_r')
// (2, 5, 'neigh_op_top_2')
// (2, 6, 'lutff_2/out')
// (2, 6, 'sp4_h_l_42')
// (2, 6, 'sp4_h_r_4')
// (2, 7, 'neigh_op_bot_2')
// (3, 5, 'neigh_op_tnl_2')
// (3, 6, 'neigh_op_lft_2')
// (3, 6, 'sp4_h_r_17')
// (3, 7, 'neigh_op_bnl_2')
// (4, 5, 'lutff_global/s_r')
// (4, 6, 'sp4_h_r_28')
// (5, 6, 'sp4_h_r_41')
// (6, 6, 'sp4_h_l_41')

reg n6 = 0;
// (0, 2, 'logic_op_tnr_2')
// (0, 3, 'logic_op_rgt_2')
// (0, 4, 'logic_op_bnr_2')
// (1, 2, 'neigh_op_top_2')
// (1, 3, 'local_g0_2')
// (1, 3, 'lutff_2/in_2')
// (1, 3, 'lutff_2/out')
// (1, 4, 'neigh_op_bot_2')
// (2, 2, 'neigh_op_tnl_2')
// (2, 3, 'local_g0_2')
// (2, 3, 'local_g1_2')
// (2, 3, 'lutff_0/in_1')
// (2, 3, 'lutff_2/in_0')
// (2, 3, 'lutff_5/in_0')
// (2, 3, 'lutff_6/in_0')
// (2, 3, 'neigh_op_lft_2')
// (2, 4, 'neigh_op_bnl_2')

reg n7 = 0;
// (0, 2, 'logic_op_tnr_3')
// (0, 3, 'logic_op_rgt_3')
// (0, 4, 'logic_op_bnr_3')
// (1, 2, 'neigh_op_top_3')
// (1, 3, 'local_g0_3')
// (1, 3, 'lutff_3/in_2')
// (1, 3, 'lutff_3/out')
// (1, 4, 'neigh_op_bot_3')
// (2, 2, 'neigh_op_tnl_3')
// (2, 3, 'local_g0_3')
// (2, 3, 'local_g1_3')
// (2, 3, 'lutff_0/in_0')
// (2, 3, 'lutff_2/in_1')
// (2, 3, 'lutff_5/in_1')
// (2, 3, 'lutff_6/in_1')
// (2, 3, 'neigh_op_lft_3')
// (2, 4, 'neigh_op_bnl_3')

reg n8 = 0;
// (0, 2, 'logic_op_tnr_4')
// (0, 3, 'logic_op_rgt_4')
// (0, 4, 'logic_op_bnr_4')
// (1, 2, 'neigh_op_top_4')
// (1, 3, 'local_g0_4')
// (1, 3, 'local_g1_4')
// (1, 3, 'lutff_1/in_2')
// (1, 3, 'lutff_4/in_2')
// (1, 3, 'lutff_4/out')
// (1, 4, 'neigh_op_bot_4')
// (2, 2, 'neigh_op_tnl_4')
// (2, 3, 'local_g0_4')
// (2, 3, 'local_g1_4')
// (2, 3, 'lutff_0/in_2')
// (2, 3, 'lutff_2/in_2')
// (2, 3, 'lutff_5/in_2')
// (2, 3, 'lutff_6/in_2')
// (2, 3, 'neigh_op_lft_4')
// (2, 4, 'neigh_op_bnl_4')

reg n9 = 0;
// (0, 2, 'span12_horz_0')
// (1, 1, 'neigh_op_tnr_6')
// (1, 1, 'sp4_r_v_b_25')
// (1, 2, 'neigh_op_rgt_6')
// (1, 2, 'sp12_h_r_3')
// (1, 2, 'sp4_r_v_b_12')
// (1, 3, 'neigh_op_bnr_6')
// (1, 3, 'sp4_r_v_b_1')
// (1, 4, 'sp4_r_v_b_41')
// (1, 5, 'sp4_r_v_b_28')
// (1, 6, 'sp4_r_v_b_17')
// (1, 7, 'sp4_r_v_b_4')
// (2, 0, 'span12_vert_15')
// (2, 0, 'span4_vert_25')
// (2, 1, 'neigh_op_top_6')
// (2, 1, 'sp12_v_b_15')
// (2, 1, 'sp4_v_b_25')
// (2, 2, 'local_g0_6')
// (2, 2, 'lutff_6/in_2')
// (2, 2, 'lutff_6/out')
// (2, 2, 'sp12_h_r_4')
// (2, 2, 'sp12_v_b_12')
// (2, 2, 'sp4_v_b_12')
// (2, 3, 'local_g1_1')
// (2, 3, 'local_g1_6')
// (2, 3, 'lutff_1/in_0')
// (2, 3, 'lutff_3/in_2')
// (2, 3, 'lutff_7/in_1')
// (2, 3, 'neigh_op_bot_6')
// (2, 3, 'sp12_v_b_11')
// (2, 3, 'sp4_v_b_1')
// (2, 3, 'sp4_v_t_41')
// (2, 4, 'sp12_v_b_8')
// (2, 4, 'sp4_v_b_41')
// (2, 5, 'sp12_v_b_7')
// (2, 5, 'sp4_v_b_28')
// (2, 6, 'local_g2_4')
// (2, 6, 'lutff_global/s_r')
// (2, 6, 'sp12_v_b_4')
// (2, 6, 'sp4_v_b_17')
// (2, 7, 'local_g0_4')
// (2, 7, 'lutff_global/s_r')
// (2, 7, 'sp12_v_b_3')
// (2, 7, 'sp4_v_b_4')
// (2, 8, 'sp12_v_b_0')
// (3, 1, 'neigh_op_tnl_6')
// (3, 2, 'neigh_op_lft_6')
// (3, 2, 'sp12_h_r_7')
// (3, 3, 'neigh_op_bnl_6')
// (4, 2, 'local_g0_0')
// (4, 2, 'lutff_5/in_1')
// (4, 2, 'sp12_h_r_8')
// (5, 2, 'sp12_h_r_11')
// (6, 2, 'sp12_h_r_12')
// (7, 2, 'sp12_h_r_15')
// (8, 2, 'sp12_h_r_16')
// (9, 2, 'sp12_h_r_19')
// (10, 2, 'sp12_h_r_20')
// (11, 2, 'sp12_h_r_23')
// (12, 2, 'sp12_h_l_23')

reg n10 = 0;
// (0, 2, 'span4_horz_0')
// (1, 1, 'neigh_op_tnr_4')
// (1, 2, 'neigh_op_rgt_4')
// (1, 2, 'sp4_h_r_13')
// (1, 2, 'sp4_r_v_b_40')
// (1, 3, 'neigh_op_bnr_4')
// (1, 3, 'sp4_r_v_b_29')
// (1, 4, 'sp4_r_v_b_16')
// (1, 5, 'sp4_r_v_b_5')
// (2, 1, 'neigh_op_top_4')
// (2, 1, 'sp4_r_v_b_36')
// (2, 1, 'sp4_v_t_40')
// (2, 2, 'local_g1_4')
// (2, 2, 'lutff_2/in_1')
// (2, 2, 'lutff_4/in_1')
// (2, 2, 'lutff_4/out')
// (2, 2, 'sp4_h_r_24')
// (2, 2, 'sp4_r_v_b_25')
// (2, 2, 'sp4_v_b_40')
// (2, 3, 'local_g2_5')
// (2, 3, 'lutff_4/in_3')
// (2, 3, 'neigh_op_bot_4')
// (2, 3, 'sp4_r_v_b_12')
// (2, 3, 'sp4_v_b_29')
// (2, 4, 'local_g1_1')
// (2, 4, 'lutff_7/in_3')
// (2, 4, 'sp4_r_v_b_1')
// (2, 4, 'sp4_v_b_16')
// (2, 5, 'sp4_h_r_5')
// (2, 5, 'sp4_v_b_5')
// (3, 0, 'span4_vert_36')
// (3, 1, 'neigh_op_tnl_4')
// (3, 1, 'sp4_v_b_36')
// (3, 2, 'neigh_op_lft_4')
// (3, 2, 'sp4_h_r_37')
// (3, 2, 'sp4_v_b_25')
// (3, 3, 'neigh_op_bnl_4')
// (3, 3, 'sp4_r_v_b_40')
// (3, 3, 'sp4_v_b_12')
// (3, 4, 'sp4_h_r_1')
// (3, 4, 'sp4_r_v_b_29')
// (3, 4, 'sp4_v_b_1')
// (3, 5, 'sp4_h_r_16')
// (3, 5, 'sp4_r_v_b_16')
// (3, 6, 'sp4_r_v_b_5')
// (4, 2, 'sp4_h_l_37')
// (4, 2, 'sp4_v_t_40')
// (4, 3, 'local_g2_0')
// (4, 3, 'lutff_0/in_2')
// (4, 3, 'sp4_v_b_40')
// (4, 4, 'sp4_h_r_12')
// (4, 4, 'sp4_v_b_29')
// (4, 5, 'sp4_h_r_29')
// (4, 5, 'sp4_v_b_16')
// (4, 6, 'sp4_v_b_5')
// (5, 2, 'sp4_r_v_b_40')
// (5, 3, 'sp4_r_v_b_29')
// (5, 4, 'local_g3_1')
// (5, 4, 'lutff_0/in_2')
// (5, 4, 'lutff_4/in_2')
// (5, 4, 'sp4_h_r_25')
// (5, 4, 'sp4_r_v_b_16')
// (5, 5, 'local_g2_0')
// (5, 5, 'local_g3_0')
// (5, 5, 'lutff_0/in_2')
// (5, 5, 'lutff_1/in_2')
// (5, 5, 'lutff_2/in_2')
// (5, 5, 'lutff_4/in_2')
// (5, 5, 'lutff_5/in_2')
// (5, 5, 'sp4_h_r_40')
// (5, 5, 'sp4_r_v_b_5')
// (6, 1, 'sp4_v_t_40')
// (6, 2, 'sp4_v_b_40')
// (6, 3, 'local_g3_5')
// (6, 3, 'lutff_2/in_2')
// (6, 3, 'lutff_4/in_2')
// (6, 3, 'sp4_v_b_29')
// (6, 4, 'local_g3_4')
// (6, 4, 'lutff_3/in_2')
// (6, 4, 'sp4_h_r_36')
// (6, 4, 'sp4_v_b_16')
// (6, 5, 'local_g0_5')
// (6, 5, 'local_g1_5')
// (6, 5, 'lutff_0/in_2')
// (6, 5, 'lutff_1/in_2')
// (6, 5, 'lutff_2/in_2')
// (6, 5, 'lutff_3/in_3')
// (6, 5, 'lutff_4/in_2')
// (6, 5, 'sp4_h_l_40')
// (6, 5, 'sp4_v_b_5')
// (7, 4, 'sp4_h_l_36')

reg n11 = 0;
// (0, 2, 'span4_horz_1')
// (0, 3, 'span12_horz_4')
// (1, 2, 'sp4_h_r_12')
// (1, 3, 'sp12_h_r_7')
// (1, 3, 'sp4_h_r_1')
// (2, 2, 'local_g3_1')
// (2, 2, 'lutff_4/in_2')
// (2, 2, 'sp4_h_r_25')
// (2, 3, 'sp12_h_r_8')
// (2, 3, 'sp4_h_r_12')
// (3, 2, 'neigh_op_tnr_2')
// (3, 2, 'sp4_h_r_36')
// (3, 3, 'neigh_op_rgt_2')
// (3, 3, 'sp12_h_r_11')
// (3, 3, 'sp4_h_r_25')
// (3, 3, 'sp4_r_v_b_36')
// (3, 4, 'neigh_op_bnr_2')
// (3, 4, 'sp4_r_v_b_25')
// (3, 5, 'sp4_h_r_1')
// (3, 5, 'sp4_r_v_b_12')
// (3, 6, 'sp4_r_v_b_1')
// (4, 0, 'span12_vert_8')
// (4, 1, 'sp12_v_b_8')
// (4, 2, 'neigh_op_top_2')
// (4, 2, 'sp12_v_b_7')
// (4, 2, 'sp4_h_l_36')
// (4, 2, 'sp4_v_t_36')
// (4, 3, 'local_g1_2')
// (4, 3, 'lutff_0/in_1')
// (4, 3, 'lutff_2/out')
// (4, 3, 'sp12_h_r_12')
// (4, 3, 'sp12_v_b_4')
// (4, 3, 'sp4_h_r_36')
// (4, 3, 'sp4_v_b_36')
// (4, 4, 'neigh_op_bot_2')
// (4, 4, 'sp12_v_b_3')
// (4, 4, 'sp4_r_v_b_36')
// (4, 4, 'sp4_v_b_25')
// (4, 5, 'sp12_h_r_0')
// (4, 5, 'sp12_v_b_0')
// (4, 5, 'sp4_h_r_12')
// (4, 5, 'sp4_r_v_b_25')
// (4, 5, 'sp4_v_b_12')
// (4, 6, 'sp4_r_v_b_12')
// (4, 6, 'sp4_v_b_1')
// (4, 7, 'sp4_r_v_b_1')
// (5, 2, 'neigh_op_tnl_2')
// (5, 3, 'neigh_op_lft_2')
// (5, 3, 'sp12_h_r_15')
// (5, 3, 'sp4_h_l_36')
// (5, 3, 'sp4_v_t_36')
// (5, 4, 'local_g3_2')
// (5, 4, 'lutff_0/in_1')
// (5, 4, 'lutff_4/in_1')
// (5, 4, 'neigh_op_bnl_2')
// (5, 4, 'sp4_v_b_36')
// (5, 5, 'local_g1_3')
// (5, 5, 'local_g2_1')
// (5, 5, 'lutff_0/in_1')
// (5, 5, 'lutff_1/in_1')
// (5, 5, 'lutff_2/in_1')
// (5, 5, 'lutff_4/in_1')
// (5, 5, 'lutff_5/in_1')
// (5, 5, 'sp12_h_r_3')
// (5, 5, 'sp4_h_r_25')
// (5, 5, 'sp4_v_b_25')
// (5, 6, 'sp4_v_b_12')
// (5, 7, 'sp4_v_b_1')
// (6, 2, 'sp4_r_v_b_36')
// (6, 3, 'local_g1_0')
// (6, 3, 'lutff_2/in_1')
// (6, 3, 'lutff_4/in_1')
// (6, 3, 'sp12_h_r_16')
// (6, 3, 'sp4_r_v_b_25')
// (6, 4, 'local_g2_4')
// (6, 4, 'lutff_3/in_1')
// (6, 4, 'sp4_r_v_b_12')
// (6, 5, 'local_g2_4')
// (6, 5, 'local_g3_4')
// (6, 5, 'lutff_0/in_1')
// (6, 5, 'lutff_1/in_1')
// (6, 5, 'lutff_2/in_1')
// (6, 5, 'lutff_3/in_2')
// (6, 5, 'lutff_4/in_1')
// (6, 5, 'sp12_h_r_4')
// (6, 5, 'sp4_h_r_36')
// (6, 5, 'sp4_r_v_b_1')
// (7, 1, 'sp4_v_t_36')
// (7, 2, 'sp4_v_b_36')
// (7, 3, 'sp12_h_r_19')
// (7, 3, 'sp4_v_b_25')
// (7, 4, 'sp4_v_b_12')
// (7, 5, 'sp12_h_r_7')
// (7, 5, 'sp4_h_l_36')
// (7, 5, 'sp4_v_b_1')
// (8, 3, 'sp12_h_r_20')
// (8, 5, 'sp12_h_r_8')
// (9, 3, 'sp12_h_r_23')
// (9, 5, 'sp12_h_r_11')
// (10, 3, 'sp12_h_l_23')
// (10, 5, 'sp12_h_r_12')
// (11, 5, 'sp12_h_r_15')
// (12, 5, 'sp12_h_r_16')
// (13, 5, 'span12_horz_16')

wire n12;
// (0, 3, 'span12_horz_0')
// (1, 2, 'neigh_op_tnr_6')
// (1, 3, 'neigh_op_rgt_6')
// (1, 3, 'sp12_h_r_3')
// (1, 4, 'neigh_op_bnr_6')
// (2, 2, 'neigh_op_top_6')
// (2, 3, 'local_g2_6')
// (2, 3, 'lutff_4/in_0')
// (2, 3, 'lutff_6/out')
// (2, 3, 'sp12_h_r_4')
// (2, 4, 'neigh_op_bot_6')
// (3, 2, 'neigh_op_tnl_6')
// (3, 3, 'neigh_op_lft_6')
// (3, 3, 'sp12_h_r_7')
// (3, 4, 'neigh_op_bnl_6')
// (4, 3, 'local_g0_0')
// (4, 3, 'local_g1_0')
// (4, 3, 'lutff_2/in_2')
// (4, 3, 'lutff_5/in_0')
// (4, 3, 'sp12_h_r_8')
// (5, 3, 'sp12_h_r_11')
// (6, 3, 'sp12_h_r_12')
// (7, 3, 'sp12_h_r_15')
// (8, 3, 'sp12_h_r_16')
// (9, 3, 'sp12_h_r_19')
// (10, 3, 'sp12_h_r_20')
// (11, 3, 'sp12_h_r_23')
// (12, 3, 'sp12_h_l_23')

reg n13 = 0;
// (0, 4, 'logic_op_tnr_2')
// (0, 5, 'logic_op_rgt_2')
// (0, 5, 'span12_horz_11')
// (0, 6, 'logic_op_bnr_2')
// (1, 3, 'sp4_r_v_b_45')
// (1, 4, 'neigh_op_top_2')
// (1, 4, 'sp4_r_v_b_32')
// (1, 5, 'local_g1_2')
// (1, 5, 'lutff_2/in_3')
// (1, 5, 'lutff_2/out')
// (1, 5, 'sp12_h_r_12')
// (1, 5, 'sp4_r_v_b_21')
// (1, 6, 'neigh_op_bot_2')
// (1, 6, 'sp4_r_v_b_8')
// (2, 2, 'sp4_v_t_45')
// (2, 3, 'sp4_v_b_45')
// (2, 4, 'neigh_op_tnl_2')
// (2, 4, 'sp4_v_b_32')
// (2, 5, 'local_g1_2')
// (2, 5, 'lutff_0/in_1')
// (2, 5, 'neigh_op_lft_2')
// (2, 5, 'sp12_h_r_15')
// (2, 5, 'sp4_v_b_21')
// (2, 6, 'local_g2_2')
// (2, 6, 'local_g3_2')
// (2, 6, 'lutff_0/in_3')
// (2, 6, 'lutff_6/in_3')
// (2, 6, 'lutff_7/in_3')
// (2, 6, 'neigh_op_bnl_2')
// (2, 6, 'sp4_h_r_8')
// (2, 6, 'sp4_v_b_8')
// (3, 5, 'sp12_h_r_16')
// (3, 6, 'sp4_h_r_21')
// (4, 5, 'local_g1_3')
// (4, 5, 'lutff_1/in_3')
// (4, 5, 'sp12_h_r_19')
// (4, 6, 'local_g2_0')
// (4, 6, 'lutff_3/in_3')
// (4, 6, 'sp4_h_r_32')
// (5, 5, 'sp12_h_r_20')
// (5, 6, 'sp4_h_r_45')
// (6, 5, 'sp12_h_r_23')
// (6, 6, 'sp4_h_l_45')
// (7, 5, 'sp12_h_l_23')

reg n14 = 0;
// (0, 4, 'span12_horz_2')
// (1, 4, 'sp12_h_r_5')
// (2, 4, 'sp12_h_r_6')
// (3, 4, 'sp12_h_r_9')
// (3, 4, 'sp4_h_r_4')
// (4, 4, 'sp12_h_r_10')
// (4, 4, 'sp4_h_r_17')
// (5, 4, 'sp12_h_r_13')
// (5, 4, 'sp4_h_r_28')
// (6, 4, 'local_g3_1')
// (6, 4, 'lutff_3/in_3')
// (6, 4, 'sp12_h_r_14')
// (6, 4, 'sp4_h_r_41')
// (7, 4, 'sp12_h_r_17')
// (7, 4, 'sp4_h_l_41')
// (8, 4, 'sp12_h_r_18')
// (9, 4, 'local_g1_5')
// (9, 4, 'lutff_0/in_0')
// (9, 4, 'sp12_h_r_21')
// (10, 4, 'neigh_op_tnr_3')
// (10, 4, 'sp12_h_r_22')
// (10, 5, 'neigh_op_rgt_3')
// (10, 6, 'neigh_op_bnr_3')
// (11, 4, 'neigh_op_top_3')
// (11, 4, 'sp12_h_l_22')
// (11, 4, 'sp12_v_t_22')
// (11, 5, 'lutff_3/out')
// (11, 5, 'sp12_v_b_22')
// (11, 6, 'neigh_op_bot_3')
// (11, 6, 'sp12_v_b_21')
// (11, 7, 'sp12_v_b_18')
// (11, 8, 'sp12_v_b_17')
// (11, 9, 'sp12_v_b_14')
// (11, 10, 'sp12_v_b_13')
// (11, 11, 'sp12_v_b_10')
// (11, 12, 'sp12_v_b_9')
// (11, 13, 'sp12_v_b_6')
// (11, 14, 'sp12_v_b_5')
// (11, 15, 'sp12_v_b_2')
// (11, 16, 'sp12_v_b_1')
// (12, 4, 'neigh_op_tnl_3')
// (12, 5, 'neigh_op_lft_3')
// (12, 6, 'neigh_op_bnl_3')

wire rst;
// (0, 4, 'span4_horz_24')
// (0, 14, 'io_1/D_IN_0')
// (0, 14, 'io_1/PAD')
// (0, 14, 'span12_horz_20')
// (1, 1, 'sp4_r_v_b_37')
// (1, 2, 'sp4_h_r_1')
// (1, 2, 'sp4_h_r_7')
// (1, 2, 'sp4_r_v_b_24')
// (1, 2, 'sp4_v_t_36')
// (1, 3, 'local_g2_4')
// (1, 3, 'lutff_global/s_r')
// (1, 3, 'sp4_r_v_b_13')
// (1, 3, 'sp4_v_b_36')
// (1, 4, 'sp4_h_r_37')
// (1, 4, 'sp4_r_v_b_0')
// (1, 4, 'sp4_v_b_25')
// (1, 5, 'sp4_r_v_b_43')
// (1, 5, 'sp4_v_b_12')
// (1, 6, 'sp4_r_v_b_30')
// (1, 6, 'sp4_v_b_1')
// (1, 7, 'sp4_r_v_b_19')
// (1, 8, 'sp4_r_v_b_6')
// (1, 13, 'neigh_op_tnl_2')
// (1, 13, 'neigh_op_tnl_6')
// (1, 14, 'neigh_op_lft_2')
// (1, 14, 'neigh_op_lft_6')
// (1, 14, 'sp12_h_r_23')
// (1, 15, 'neigh_op_bnl_2')
// (1, 15, 'neigh_op_bnl_6')
// (2, 0, 'span4_vert_37')
// (2, 1, 'sp4_v_b_37')
// (2, 2, 'local_g1_0')
// (2, 2, 'lutff_2/in_3')
// (2, 2, 'lutff_4/in_3')
// (2, 2, 'lutff_6/in_3')
// (2, 2, 'sp12_h_r_0')
// (2, 2, 'sp12_v_t_23')
// (2, 2, 'sp4_h_r_12')
// (2, 2, 'sp4_h_r_18')
// (2, 2, 'sp4_v_b_24')
// (2, 3, 'local_g1_5')
// (2, 3, 'local_g3_7')
// (2, 3, 'lutff_3/in_1')
// (2, 3, 'lutff_global/s_r')
// (2, 3, 'sp12_v_b_23')
// (2, 3, 'sp4_v_b_13')
// (2, 4, 'sp12_v_b_20')
// (2, 4, 'sp4_h_l_37')
// (2, 4, 'sp4_v_b_0')
// (2, 4, 'sp4_v_t_43')
// (2, 5, 'sp12_v_b_19')
// (2, 5, 'sp4_v_b_43')
// (2, 6, 'local_g2_6')
// (2, 6, 'local_g3_0')
// (2, 6, 'lutff_1/in_3')
// (2, 6, 'lutff_2/in_3')
// (2, 6, 'sp12_v_b_16')
// (2, 6, 'sp4_v_b_30')
// (2, 7, 'sp12_v_b_15')
// (2, 7, 'sp4_v_b_19')
// (2, 8, 'local_g2_4')
// (2, 8, 'lutff_3/in_3')
// (2, 8, 'sp12_v_b_12')
// (2, 8, 'sp4_v_b_6')
// (2, 9, 'sp12_v_b_11')
// (2, 10, 'sp12_v_b_8')
// (2, 11, 'sp12_v_b_7')
// (2, 12, 'sp12_v_b_4')
// (2, 13, 'sp12_v_b_3')
// (2, 14, 'sp12_h_l_23')
// (2, 14, 'sp12_v_b_0')
// (3, 2, 'sp12_h_r_3')
// (3, 2, 'sp4_h_r_25')
// (3, 2, 'sp4_h_r_31')
// (4, 2, 'local_g0_4')
// (4, 2, 'lutff_7/in_3')
// (4, 2, 'sp12_h_r_4')
// (4, 2, 'sp4_h_r_36')
// (4, 2, 'sp4_h_r_42')
// (4, 3, 'local_g2_4')
// (4, 3, 'local_g2_5')
// (4, 3, 'lutff_2/in_1')
// (4, 3, 'lutff_5/in_3')
// (4, 3, 'sp4_r_v_b_36')
// (4, 3, 'sp4_r_v_b_37')
// (4, 4, 'sp4_r_v_b_24')
// (4, 4, 'sp4_r_v_b_25')
// (4, 5, 'sp4_r_v_b_12')
// (4, 5, 'sp4_r_v_b_13')
// (4, 6, 'sp4_r_v_b_0')
// (4, 6, 'sp4_r_v_b_1')
// (5, 2, 'sp12_h_r_7')
// (5, 2, 'sp4_h_l_36')
// (5, 2, 'sp4_h_l_42')
// (5, 2, 'sp4_v_t_36')
// (5, 2, 'sp4_v_t_37')
// (5, 3, 'sp4_v_b_36')
// (5, 3, 'sp4_v_b_37')
// (5, 4, 'sp4_v_b_24')
// (5, 4, 'sp4_v_b_25')
// (5, 5, 'sp4_v_b_12')
// (5, 5, 'sp4_v_b_13')
// (5, 6, 'sp4_v_b_0')
// (5, 6, 'sp4_v_b_1')
// (6, 2, 'sp12_h_r_8')
// (7, 2, 'sp12_h_r_11')
// (8, 2, 'sp12_h_r_12')
// (9, 2, 'sp12_h_r_15')
// (10, 2, 'sp12_h_r_16')
// (11, 2, 'sp12_h_r_19')
// (12, 2, 'sp12_h_r_20')
// (13, 2, 'span12_horz_20')

reg n16 = 0;
// (0, 5, 'logic_op_tnr_6')
// (0, 6, 'logic_op_rgt_6')
// (0, 6, 'span12_horz_3')
// (0, 7, 'logic_op_bnr_6')
// (1, 5, 'neigh_op_top_6')
// (1, 6, 'lutff_6/out')
// (1, 6, 'sp12_h_r_4')
// (1, 6, 'sp4_r_v_b_45')
// (1, 7, 'neigh_op_bot_6')
// (1, 7, 'sp4_r_v_b_32')
// (1, 8, 'sp4_r_v_b_21')
// (1, 9, 'sp4_r_v_b_8')
// (2, 5, 'neigh_op_tnl_6')
// (2, 5, 'sp4_h_r_8')
// (2, 5, 'sp4_v_t_45')
// (2, 6, 'neigh_op_lft_6')
// (2, 6, 'sp12_h_r_7')
// (2, 6, 'sp4_v_b_45')
// (2, 7, 'neigh_op_bnl_6')
// (2, 7, 'sp4_v_b_32')
// (2, 8, 'sp4_v_b_21')
// (2, 9, 'sp4_v_b_8')
// (3, 5, 'sp4_h_r_21')
// (3, 6, 'sp12_h_r_8')
// (4, 5, 'sp4_h_r_32')
// (4, 6, 'sp12_h_r_11')
// (5, 5, 'local_g2_5')
// (5, 5, 'lutff_0/in_3')
// (5, 5, 'sp4_h_r_45')
// (5, 6, 'local_g0_4')
// (5, 6, 'lutff_6/in_0')
// (5, 6, 'sp12_h_r_12')
// (6, 5, 'sp4_h_l_45')
// (6, 6, 'sp12_h_r_15')
// (7, 6, 'sp12_h_r_16')
// (8, 6, 'sp12_h_r_19')
// (9, 6, 'sp12_h_r_20')
// (10, 6, 'sp12_h_r_23')
// (11, 6, 'sp12_h_l_23')

reg n17 = 0;
// (0, 5, 'logic_op_tnr_7')
// (0, 6, 'logic_op_rgt_7')
// (0, 7, 'logic_op_bnr_7')
// (1, 5, 'neigh_op_top_7')
// (1, 6, 'local_g1_7')
// (1, 6, 'lutff_6/in_0')
// (1, 6, 'lutff_7/out')
// (1, 7, 'neigh_op_bot_7')
// (2, 5, 'neigh_op_tnl_7')
// (2, 6, 'neigh_op_lft_7')
// (2, 7, 'neigh_op_bnl_7')

wire n18;
// (0, 5, 'span12_horz_0')
// (1, 5, 'sp12_h_r_3')
// (1, 6, 'sp4_h_r_9')
// (2, 5, 'sp12_h_r_4')
// (2, 6, 'local_g0_4')
// (2, 6, 'lutff_5/in_1')
// (2, 6, 'sp4_h_r_20')
// (3, 4, 'neigh_op_tnr_0')
// (3, 5, 'neigh_op_rgt_0')
// (3, 5, 'sp12_h_r_7')
// (3, 6, 'neigh_op_bnr_0')
// (3, 6, 'sp4_h_r_33')
// (4, 3, 'sp4_r_v_b_41')
// (4, 4, 'neigh_op_top_0')
// (4, 4, 'sp4_r_v_b_28')
// (4, 5, 'lutff_0/out')
// (4, 5, 'sp12_h_r_8')
// (4, 5, 'sp4_r_v_b_17')
// (4, 6, 'neigh_op_bot_0')
// (4, 6, 'sp4_h_r_44')
// (4, 6, 'sp4_r_v_b_4')
// (5, 2, 'sp4_v_t_41')
// (5, 3, 'sp4_v_b_41')
// (5, 4, 'neigh_op_tnl_0')
// (5, 4, 'sp4_v_b_28')
// (5, 5, 'neigh_op_lft_0')
// (5, 5, 'sp12_h_r_11')
// (5, 5, 'sp4_v_b_17')
// (5, 6, 'neigh_op_bnl_0')
// (5, 6, 'sp4_h_l_44')
// (5, 6, 'sp4_v_b_4')
// (6, 5, 'sp12_h_r_12')
// (7, 5, 'local_g0_7')
// (7, 5, 'lutff_7/in_2')
// (7, 5, 'sp12_h_r_15')
// (8, 5, 'local_g0_0')
// (8, 5, 'lutff_3/in_1')
// (8, 5, 'sp12_h_r_16')
// (9, 5, 'sp12_h_r_19')
// (10, 5, 'sp12_h_r_20')
// (11, 5, 'sp12_h_r_23')
// (12, 5, 'sp12_h_l_23')

reg n19 = 0;
// (0, 5, 'span12_horz_14')
// (1, 4, 'neigh_op_tnr_5')
// (1, 5, 'neigh_op_rgt_5')
// (1, 5, 'sp12_h_r_1')
// (1, 5, 'sp12_h_r_17')
// (1, 6, 'neigh_op_bnr_5')
// (2, 4, 'neigh_op_top_5')
// (2, 5, 'local_g0_5')
// (2, 5, 'lutff_5/in_2')
// (2, 5, 'lutff_5/out')
// (2, 5, 'sp12_h_r_18')
// (2, 5, 'sp12_h_r_2')
// (2, 5, 'sp4_r_v_b_43')
// (2, 6, 'local_g0_6')
// (2, 6, 'lutff_3/in_3')
// (2, 6, 'neigh_op_bot_5')
// (2, 6, 'sp4_r_v_b_30')
// (2, 7, 'sp4_r_v_b_19')
// (2, 8, 'sp4_r_v_b_6')
// (3, 4, 'neigh_op_tnl_5')
// (3, 4, 'sp4_v_t_43')
// (3, 5, 'neigh_op_lft_5')
// (3, 5, 'sp12_h_r_21')
// (3, 5, 'sp12_h_r_5')
// (3, 5, 'sp4_v_b_43')
// (3, 6, 'neigh_op_bnl_5')
// (3, 6, 'sp4_v_b_30')
// (3, 7, 'sp4_v_b_19')
// (3, 8, 'sp4_v_b_6')
// (4, 5, 'local_g1_6')
// (4, 5, 'lutff_0/in_3')
// (4, 5, 'sp12_h_r_22')
// (4, 5, 'sp12_h_r_6')
// (4, 5, 'sp4_r_v_b_46')
// (4, 6, 'local_g2_3')
// (4, 6, 'lutff_0/in_1')
// (4, 6, 'lutff_4/in_1')
// (4, 6, 'sp4_r_v_b_35')
// (4, 7, 'sp4_r_v_b_22')
// (4, 7, 'sp4_r_v_b_44')
// (4, 8, 'sp4_r_v_b_11')
// (4, 8, 'sp4_r_v_b_33')
// (4, 9, 'sp4_r_v_b_20')
// (4, 10, 'sp4_r_v_b_9')
// (5, 4, 'sp4_v_t_46')
// (5, 5, 'sp12_h_l_22')
// (5, 5, 'sp12_h_r_9')
// (5, 5, 'sp12_v_t_22')
// (5, 5, 'sp4_v_b_46')
// (5, 6, 'sp12_v_b_22')
// (5, 6, 'sp4_h_r_9')
// (5, 6, 'sp4_v_b_35')
// (5, 6, 'sp4_v_t_44')
// (5, 7, 'sp12_v_b_21')
// (5, 7, 'sp4_v_b_22')
// (5, 7, 'sp4_v_b_44')
// (5, 8, 'sp12_v_b_18')
// (5, 8, 'sp4_v_b_11')
// (5, 8, 'sp4_v_b_33')
// (5, 9, 'sp12_v_b_17')
// (5, 9, 'sp4_v_b_20')
// (5, 10, 'sp12_v_b_14')
// (5, 10, 'sp4_v_b_9')
// (5, 11, 'sp12_v_b_13')
// (5, 12, 'sp12_v_b_10')
// (5, 13, 'sp12_v_b_9')
// (5, 14, 'sp12_v_b_6')
// (5, 15, 'sp12_v_b_5')
// (5, 16, 'sp12_v_b_2')
// (5, 17, 'span12_vert_1')
// (6, 5, 'sp12_h_r_10')
// (6, 6, 'sp4_h_r_20')
// (7, 5, 'local_g1_5')
// (7, 5, 'lutff_2/in_2')
// (7, 5, 'lutff_5/in_1')
// (7, 5, 'sp12_h_r_13')
// (7, 6, 'local_g2_1')
// (7, 6, 'lutff_3/in_2')
// (7, 6, 'lutff_4/in_1')
// (7, 6, 'sp4_h_r_33')
// (8, 5, 'sp12_h_r_14')
// (8, 6, 'sp4_h_r_44')
// (9, 5, 'sp12_h_r_17')
// (9, 6, 'sp4_h_l_44')
// (10, 5, 'sp12_h_r_18')
// (11, 5, 'sp12_h_r_21')
// (12, 5, 'sp12_h_r_22')
// (13, 5, 'span12_horz_22')

reg n20 = 0;
// (0, 5, 'span12_horz_2')
// (0, 6, 'span4_horz_0')
// (1, 5, 'sp12_h_r_5')
// (1, 6, 'sp4_h_r_13')
// (2, 5, 'local_g1_6')
// (2, 5, 'lutff_1/in_2')
// (2, 5, 'sp12_h_r_6')
// (2, 6, 'local_g2_0')
// (2, 6, 'lutff_0/in_0')
// (2, 6, 'lutff_6/in_2')
// (2, 6, 'lutff_7/in_1')
// (2, 6, 'sp4_h_r_24')
// (3, 3, 'sp4_r_v_b_42')
// (3, 4, 'neigh_op_tnr_1')
// (3, 4, 'sp4_r_v_b_31')
// (3, 5, 'neigh_op_rgt_1')
// (3, 5, 'sp12_h_r_9')
// (3, 5, 'sp4_r_v_b_18')
// (3, 6, 'neigh_op_bnr_1')
// (3, 6, 'sp4_h_r_37')
// (3, 6, 'sp4_r_v_b_7')
// (4, 2, 'sp4_v_t_42')
// (4, 3, 'sp4_v_b_42')
// (4, 4, 'neigh_op_top_1')
// (4, 4, 'sp4_v_b_31')
// (4, 5, 'local_g0_1')
// (4, 5, 'lutff_1/in_2')
// (4, 5, 'lutff_1/out')
// (4, 5, 'sp12_h_r_10')
// (4, 5, 'sp4_v_b_18')
// (4, 6, 'local_g0_7')
// (4, 6, 'lutff_3/in_2')
// (4, 6, 'neigh_op_bot_1')
// (4, 6, 'sp4_h_l_37')
// (4, 6, 'sp4_v_b_7')
// (5, 4, 'neigh_op_tnl_1')
// (5, 5, 'neigh_op_lft_1')
// (5, 5, 'sp12_h_r_13')
// (5, 6, 'neigh_op_bnl_1')
// (6, 5, 'sp12_h_r_14')
// (7, 5, 'sp12_h_r_17')
// (8, 5, 'sp12_h_r_18')
// (9, 5, 'sp12_h_r_21')
// (10, 5, 'sp12_h_r_22')
// (11, 5, 'sp12_h_l_22')

reg n21 = 0;
// (0, 5, 'span4_horz_20')
// (0, 5, 'span4_horz_4')
// (1, 4, 'neigh_op_tnr_6')
// (1, 5, 'neigh_op_rgt_6')
// (1, 5, 'sp4_h_r_17')
// (1, 5, 'sp4_h_r_33')
// (1, 6, 'neigh_op_bnr_6')
// (2, 3, 'sp4_r_v_b_37')
// (2, 4, 'neigh_op_top_6')
// (2, 4, 'sp4_r_v_b_24')
// (2, 5, 'local_g0_6')
// (2, 5, 'lutff_6/in_2')
// (2, 5, 'lutff_6/out')
// (2, 5, 'sp4_h_r_28')
// (2, 5, 'sp4_h_r_44')
// (2, 5, 'sp4_r_v_b_13')
// (2, 6, 'local_g1_6')
// (2, 6, 'lutff_3/in_0')
// (2, 6, 'neigh_op_bot_6')
// (2, 6, 'sp4_r_v_b_0')
// (3, 2, 'sp4_v_t_37')
// (3, 3, 'sp4_v_b_37')
// (3, 4, 'neigh_op_tnl_6')
// (3, 4, 'sp4_v_b_24')
// (3, 5, 'neigh_op_lft_6')
// (3, 5, 'sp4_h_l_44')
// (3, 5, 'sp4_h_r_41')
// (3, 5, 'sp4_h_r_5')
// (3, 5, 'sp4_v_b_13')
// (3, 6, 'neigh_op_bnl_6')
// (3, 6, 'sp4_h_r_0')
// (3, 6, 'sp4_v_b_0')
// (4, 5, 'local_g0_0')
// (4, 5, 'lutff_0/in_2')
// (4, 5, 'sp4_h_l_41')
// (4, 5, 'sp4_h_r_16')
// (4, 5, 'sp4_h_r_4')
// (4, 6, 'local_g1_5')
// (4, 6, 'lutff_1/in_3')
// (4, 6, 'sp4_h_r_13')
// (5, 5, 'sp4_h_r_17')
// (5, 5, 'sp4_h_r_29')
// (5, 6, 'sp4_h_r_24')
// (6, 5, 'sp4_h_r_28')
// (6, 5, 'sp4_h_r_40')
// (6, 6, 'sp4_h_r_37')
// (6, 6, 'sp4_r_v_b_40')
// (6, 7, 'sp4_r_v_b_29')
// (6, 8, 'sp4_r_v_b_16')
// (6, 9, 'sp4_r_v_b_5')
// (7, 5, 'local_g0_0')
// (7, 5, 'local_g2_1')
// (7, 5, 'lutff_0/in_2')
// (7, 5, 'lutff_5/in_2')
// (7, 5, 'sp4_h_l_40')
// (7, 5, 'sp4_h_r_41')
// (7, 5, 'sp4_h_r_8')
// (7, 5, 'sp4_v_t_40')
// (7, 6, 'local_g2_0')
// (7, 6, 'lutff_4/in_0')
// (7, 6, 'lutff_6/in_0')
// (7, 6, 'sp4_h_l_37')
// (7, 6, 'sp4_v_b_40')
// (7, 7, 'sp4_v_b_29')
// (7, 8, 'sp4_v_b_16')
// (7, 9, 'sp4_v_b_5')
// (8, 5, 'sp4_h_l_41')
// (8, 5, 'sp4_h_r_21')
// (9, 5, 'sp4_h_r_32')
// (10, 5, 'sp4_h_r_45')
// (11, 5, 'sp4_h_l_45')

reg n22 = 0;
// (0, 5, 'span4_horz_6')
// (1, 3, 'sp4_r_v_b_38')
// (1, 4, 'neigh_op_tnr_7')
// (1, 4, 'sp4_r_v_b_27')
// (1, 5, 'neigh_op_rgt_7')
// (1, 5, 'sp4_h_r_19')
// (1, 5, 'sp4_r_v_b_14')
// (1, 6, 'neigh_op_bnr_7')
// (1, 6, 'sp4_r_v_b_3')
// (2, 2, 'sp4_v_t_38')
// (2, 3, 'sp4_v_b_38')
// (2, 4, 'neigh_op_top_7')
// (2, 4, 'sp4_v_b_27')
// (2, 5, 'local_g0_7')
// (2, 5, 'lutff_7/in_2')
// (2, 5, 'lutff_7/out')
// (2, 5, 'sp4_h_r_30')
// (2, 5, 'sp4_v_b_14')
// (2, 6, 'local_g0_7')
// (2, 6, 'lutff_3/in_2')
// (2, 6, 'lutff_5/in_2')
// (2, 6, 'neigh_op_bot_7')
// (2, 6, 'sp4_h_r_9')
// (2, 6, 'sp4_v_b_3')
// (3, 4, 'neigh_op_tnl_7')
// (3, 5, 'neigh_op_lft_7')
// (3, 5, 'sp4_h_r_43')
// (3, 6, 'neigh_op_bnl_7')
// (3, 6, 'sp4_h_r_20')
// (4, 5, 'sp4_h_l_43')
// (4, 5, 'sp4_h_r_6')
// (4, 6, 'local_g2_1')
// (4, 6, 'lutff_1/in_2')
// (4, 6, 'sp4_h_r_33')
// (5, 5, 'sp4_h_r_19')
// (5, 6, 'sp4_h_r_44')
// (5, 7, 'sp4_r_v_b_39')
// (5, 8, 'sp4_r_v_b_26')
// (5, 9, 'sp4_r_v_b_15')
// (5, 10, 'sp4_r_v_b_2')
// (6, 5, 'sp4_h_r_30')
// (6, 6, 'sp4_h_l_44')
// (6, 6, 'sp4_h_r_5')
// (6, 6, 'sp4_h_r_7')
// (6, 6, 'sp4_v_t_39')
// (6, 7, 'sp4_v_b_39')
// (6, 8, 'sp4_v_b_26')
// (6, 9, 'sp4_v_b_15')
// (6, 10, 'sp4_v_b_2')
// (7, 5, 'local_g2_3')
// (7, 5, 'local_g3_3')
// (7, 5, 'lutff_0/in_1')
// (7, 5, 'lutff_4/in_2')
// (7, 5, 'lutff_5/in_0')
// (7, 5, 'lutff_7/in_0')
// (7, 5, 'sp4_h_r_43')
// (7, 6, 'local_g0_0')
// (7, 6, 'local_g1_2')
// (7, 6, 'lutff_4/in_2')
// (7, 6, 'lutff_6/in_1')
// (7, 6, 'sp4_h_r_16')
// (7, 6, 'sp4_h_r_18')
// (8, 5, 'sp4_h_l_43')
// (8, 6, 'sp4_h_r_29')
// (8, 6, 'sp4_h_r_31')
// (9, 6, 'sp4_h_r_40')
// (9, 6, 'sp4_h_r_42')
// (10, 6, 'sp4_h_l_40')
// (10, 6, 'sp4_h_l_42')

reg n23 = 0;
// (0, 6, 'logic_op_tnr_4')
// (0, 7, 'logic_op_rgt_4')
// (0, 8, 'logic_op_bnr_4')
// (1, 6, 'local_g1_4')
// (1, 6, 'lutff_7/in_0')
// (1, 6, 'neigh_op_top_4')
// (1, 7, 'lutff_4/out')
// (1, 8, 'neigh_op_bot_4')
// (2, 6, 'neigh_op_tnl_4')
// (2, 7, 'neigh_op_lft_4')
// (2, 8, 'neigh_op_bnl_4')

reg n24 = 0;
// (0, 6, 'span4_horz_1')
// (0, 6, 'span4_horz_25')
// (1, 6, 'sp4_h_r_12')
// (1, 6, 'sp4_h_r_36')
// (2, 6, 'sp4_h_l_36')
// (2, 6, 'sp4_h_r_1')
// (2, 6, 'sp4_h_r_25')
// (3, 6, 'sp12_h_r_0')
// (3, 6, 'sp4_h_r_12')
// (3, 6, 'sp4_h_r_36')
// (3, 7, 'sp4_r_v_b_43')
// (3, 8, 'sp4_r_v_b_30')
// (3, 9, 'sp4_r_v_b_19')
// (3, 10, 'sp4_r_v_b_6')
// (4, 6, 'sp12_h_r_3')
// (4, 6, 'sp4_h_l_36')
// (4, 6, 'sp4_h_r_25')
// (4, 6, 'sp4_v_t_43')
// (4, 7, 'sp4_v_b_43')
// (4, 8, 'sp4_v_b_30')
// (4, 9, 'local_g0_3')
// (4, 9, 'lutff_1/in_0')
// (4, 9, 'sp4_v_b_19')
// (4, 10, 'sp4_v_b_6')
// (5, 6, 'sp12_h_r_4')
// (5, 6, 'sp4_h_r_36')
// (5, 7, 'sp4_r_v_b_43')
// (5, 8, 'sp4_r_v_b_30')
// (5, 9, 'sp4_r_v_b_19')
// (5, 10, 'sp4_r_v_b_6')
// (6, 6, 'sp12_h_r_7')
// (6, 6, 'sp4_h_l_36')
// (6, 6, 'sp4_v_t_43')
// (6, 7, 'sp4_v_b_43')
// (6, 8, 'sp4_v_b_30')
// (6, 9, 'local_g0_3')
// (6, 9, 'lutff_3/in_2')
// (6, 9, 'lutff_7/in_2')
// (6, 9, 'sp4_v_b_19')
// (6, 10, 'sp4_v_b_6')
// (7, 6, 'local_g1_0')
// (7, 6, 'lutff_7/in_0')
// (7, 6, 'sp12_h_r_8')
// (8, 6, 'sp12_h_r_11')
// (9, 6, 'sp12_h_r_12')
// (10, 5, 'neigh_op_tnr_4')
// (10, 6, 'neigh_op_rgt_4')
// (10, 6, 'sp12_h_r_15')
// (10, 7, 'neigh_op_bnr_4')
// (11, 5, 'neigh_op_top_4')
// (11, 6, 'lutff_4/out')
// (11, 6, 'sp12_h_r_16')
// (11, 7, 'neigh_op_bot_4')
// (12, 5, 'neigh_op_tnl_4')
// (12, 6, 'neigh_op_lft_4')
// (12, 6, 'sp12_h_r_19')
// (12, 7, 'neigh_op_bnl_4')
// (13, 6, 'span12_horz_19')

reg n25 = 0;
// (0, 6, 'span4_horz_4')
// (1, 5, 'neigh_op_tnr_6')
// (1, 6, 'neigh_op_rgt_6')
// (1, 6, 'sp4_h_r_1')
// (1, 6, 'sp4_h_r_17')
// (1, 7, 'neigh_op_bnr_6')
// (2, 0, 'span12_vert_23')
// (2, 1, 'sp12_v_b_23')
// (2, 2, 'sp12_v_b_20')
// (2, 3, 'sp12_v_b_19')
// (2, 4, 'sp12_v_b_16')
// (2, 5, 'neigh_op_top_6')
// (2, 5, 'sp12_v_b_15')
// (2, 6, 'lutff_6/out')
// (2, 6, 'sp12_v_b_12')
// (2, 6, 'sp4_h_r_12')
// (2, 6, 'sp4_h_r_28')
// (2, 6, 'sp4_r_v_b_45')
// (2, 7, 'neigh_op_bot_6')
// (2, 7, 'sp12_v_b_11')
// (2, 7, 'sp4_r_v_b_32')
// (2, 8, 'sp12_v_b_8')
// (2, 8, 'sp4_r_v_b_21')
// (2, 9, 'sp12_v_b_7')
// (2, 9, 'sp4_r_v_b_8')
// (2, 10, 'sp12_v_b_4')
// (2, 11, 'sp12_v_b_3')
// (2, 12, 'sp12_h_r_0')
// (2, 12, 'sp12_v_b_0')
// (3, 5, 'neigh_op_tnl_6')
// (3, 5, 'sp4_v_t_45')
// (3, 6, 'neigh_op_lft_6')
// (3, 6, 'sp4_h_r_25')
// (3, 6, 'sp4_h_r_41')
// (3, 6, 'sp4_v_b_45')
// (3, 7, 'neigh_op_bnl_6')
// (3, 7, 'sp4_r_v_b_44')
// (3, 7, 'sp4_v_b_32')
// (3, 8, 'sp4_r_v_b_33')
// (3, 8, 'sp4_v_b_21')
// (3, 9, 'sp4_h_r_8')
// (3, 9, 'sp4_r_v_b_20')
// (3, 9, 'sp4_v_b_8')
// (3, 10, 'sp4_r_v_b_9')
// (3, 12, 'sp12_h_r_3')
// (4, 6, 'sp4_h_l_41')
// (4, 6, 'sp4_h_r_36')
// (4, 6, 'sp4_v_t_44')
// (4, 7, 'sp4_r_v_b_43')
// (4, 7, 'sp4_v_b_44')
// (4, 8, 'sp4_r_v_b_30')
// (4, 8, 'sp4_v_b_33')
// (4, 9, 'local_g0_4')
// (4, 9, 'lutff_3/in_3')
// (4, 9, 'sp4_h_r_21')
// (4, 9, 'sp4_r_v_b_19')
// (4, 9, 'sp4_v_b_20')
// (4, 10, 'sp4_h_r_9')
// (4, 10, 'sp4_r_v_b_6')
// (4, 10, 'sp4_v_b_9')
// (4, 11, 'sp4_r_v_b_43')
// (4, 12, 'sp12_h_r_4')
// (4, 12, 'sp4_r_v_b_30')
// (4, 13, 'sp4_r_v_b_19')
// (4, 14, 'sp4_h_r_8')
// (4, 14, 'sp4_r_v_b_6')
// (5, 6, 'sp4_h_l_36')
// (5, 6, 'sp4_v_t_43')
// (5, 7, 'sp4_v_b_43')
// (5, 8, 'sp4_v_b_30')
// (5, 9, 'local_g0_3')
// (5, 9, 'lutff_7/in_2')
// (5, 9, 'sp4_h_r_32')
// (5, 9, 'sp4_v_b_19')
// (5, 10, 'local_g1_4')
// (5, 10, 'lutff_1/in_2')
// (5, 10, 'sp4_h_r_20')
// (5, 10, 'sp4_v_b_6')
// (5, 10, 'sp4_v_t_43')
// (5, 11, 'local_g2_3')
// (5, 11, 'local_g3_3')
// (5, 11, 'lutff_0/in_3')
// (5, 11, 'lutff_5/in_2')
// (5, 11, 'lutff_7/in_3')
// (5, 11, 'sp4_v_b_43')
// (5, 12, 'sp12_h_r_7')
// (5, 12, 'sp4_v_b_30')
// (5, 13, 'local_g0_3')
// (5, 13, 'local_g1_3')
// (5, 13, 'lutff_0/in_3')
// (5, 13, 'lutff_1/in_3')
// (5, 13, 'lutff_2/in_2')
// (5, 13, 'sp4_v_b_19')
// (5, 14, 'local_g0_5')
// (5, 14, 'local_g1_5')
// (5, 14, 'lutff_4/in_3')
// (5, 14, 'lutff_6/in_2')
// (5, 14, 'sp4_h_r_21')
// (5, 14, 'sp4_v_b_6')
// (6, 9, 'local_g2_5')
// (6, 9, 'local_g3_5')
// (6, 9, 'lutff_2/in_3')
// (6, 9, 'lutff_4/in_2')
// (6, 9, 'sp4_h_r_45')
// (6, 10, 'sp4_h_r_33')
// (6, 10, 'sp4_r_v_b_45')
// (6, 11, 'local_g0_3')
// (6, 11, 'lutff_2/in_3')
// (6, 11, 'sp4_r_v_b_32')
// (6, 12, 'local_g1_0')
// (6, 12, 'local_g3_5')
// (6, 12, 'lutff_0/in_2')
// (6, 12, 'lutff_2/in_3')
// (6, 12, 'lutff_3/in_2')
// (6, 12, 'lutff_6/in_2')
// (6, 12, 'sp12_h_r_8')
// (6, 12, 'sp4_r_v_b_21')
// (6, 13, 'local_g2_0')
// (6, 13, 'lutff_6/in_2')
// (6, 13, 'lutff_7/in_3')
// (6, 13, 'sp4_r_v_b_8')
// (6, 14, 'sp4_h_r_32')
// (7, 7, 'sp4_r_v_b_38')
// (7, 7, 'sp4_r_v_b_44')
// (7, 8, 'sp4_r_v_b_27')
// (7, 8, 'sp4_r_v_b_33')
// (7, 9, 'sp4_h_l_45')
// (7, 9, 'sp4_r_v_b_14')
// (7, 9, 'sp4_r_v_b_20')
// (7, 9, 'sp4_v_t_45')
// (7, 10, 'local_g1_3')
// (7, 10, 'local_g2_1')
// (7, 10, 'lutff_2/in_2')
// (7, 10, 'lutff_3/in_3')
// (7, 10, 'lutff_7/in_2')
// (7, 10, 'sp4_h_r_44')
// (7, 10, 'sp4_r_v_b_3')
// (7, 10, 'sp4_r_v_b_9')
// (7, 10, 'sp4_v_b_45')
// (7, 11, 'local_g2_6')
// (7, 11, 'lutff_2/in_2')
// (7, 11, 'sp4_r_v_b_38')
// (7, 11, 'sp4_v_b_32')
// (7, 12, 'local_g0_3')
// (7, 12, 'lutff_2/in_3')
// (7, 12, 'sp12_h_r_11')
// (7, 12, 'sp4_r_v_b_27')
// (7, 12, 'sp4_v_b_21')
// (7, 13, 'local_g2_6')
// (7, 13, 'lutff_3/in_3')
// (7, 13, 'sp4_r_v_b_14')
// (7, 13, 'sp4_v_b_8')
// (7, 14, 'local_g2_5')
// (7, 14, 'lutff_0/in_3')
// (7, 14, 'lutff_1/in_2')
// (7, 14, 'lutff_2/in_3')
// (7, 14, 'lutff_5/in_2')
// (7, 14, 'sp4_h_r_45')
// (7, 14, 'sp4_r_v_b_3')
// (8, 6, 'sp4_v_t_38')
// (8, 6, 'sp4_v_t_44')
// (8, 7, 'sp4_v_b_38')
// (8, 7, 'sp4_v_b_44')
// (8, 8, 'sp4_v_b_27')
// (8, 8, 'sp4_v_b_33')
// (8, 9, 'sp4_v_b_14')
// (8, 9, 'sp4_v_b_20')
// (8, 10, 'sp4_h_l_44')
// (8, 10, 'sp4_v_b_3')
// (8, 10, 'sp4_v_b_9')
// (8, 10, 'sp4_v_t_38')
// (8, 11, 'local_g2_6')
// (8, 11, 'local_g3_6')
// (8, 11, 'lutff_0/in_3')
// (8, 11, 'lutff_7/in_3')
// (8, 11, 'sp4_v_b_38')
// (8, 12, 'local_g3_3')
// (8, 12, 'lutff_2/in_2')
// (8, 12, 'sp12_h_r_12')
// (8, 12, 'sp4_v_b_27')
// (8, 13, 'sp4_v_b_14')
// (8, 14, 'sp4_h_l_45')
// (8, 14, 'sp4_v_b_3')
// (9, 12, 'sp12_h_r_15')
// (10, 12, 'sp12_h_r_16')
// (11, 12, 'sp12_h_r_19')
// (12, 12, 'sp12_h_r_20')
// (13, 12, 'span12_horz_20')

wire select;
// (0, 7, 'span12_horz_0')
// (1, 7, 'sp12_h_r_3')
// (2, 7, 'sp12_h_r_4')
// (3, 4, 'sp4_r_v_b_40')
// (3, 5, 'sp4_r_v_b_29')
// (3, 6, 'sp4_r_v_b_16')
// (3, 7, 'sp12_h_r_7')
// (3, 7, 'sp4_r_v_b_5')
// (4, 3, 'sp4_v_t_40')
// (4, 4, 'sp4_r_v_b_42')
// (4, 4, 'sp4_v_b_40')
// (4, 5, 'sp4_r_v_b_31')
// (4, 5, 'sp4_v_b_29')
// (4, 6, 'local_g1_0')
// (4, 6, 'lutff_6/in_3')
// (4, 6, 'sp4_r_v_b_18')
// (4, 6, 'sp4_v_b_16')
// (4, 7, 'sp12_h_r_8')
// (4, 7, 'sp4_h_r_5')
// (4, 7, 'sp4_r_v_b_7')
// (4, 7, 'sp4_v_b_5')
// (5, 3, 'sp4_v_t_42')
// (5, 4, 'sp4_v_b_42')
// (5, 5, 'sp4_v_b_31')
// (5, 6, 'local_g1_2')
// (5, 6, 'lutff_2/in_3')
// (5, 6, 'sp4_v_b_18')
// (5, 7, 'sp12_h_r_11')
// (5, 7, 'sp4_h_r_16')
// (5, 7, 'sp4_h_r_7')
// (5, 7, 'sp4_v_b_7')
// (6, 7, 'sp12_h_r_12')
// (6, 7, 'sp4_h_r_18')
// (6, 7, 'sp4_h_r_29')
// (7, 7, 'sp12_h_r_15')
// (7, 7, 'sp4_h_r_31')
// (7, 7, 'sp4_h_r_40')
// (8, 7, 'sp12_h_r_16')
// (8, 7, 'sp4_h_l_40')
// (8, 7, 'sp4_h_r_2')
// (8, 7, 'sp4_h_r_42')
// (9, 7, 'sp12_h_r_19')
// (9, 7, 'sp4_h_l_42')
// (9, 7, 'sp4_h_r_15')
// (10, 7, 'sp12_h_r_20')
// (10, 7, 'sp4_h_r_26')
// (11, 6, 'local_g2_7')
// (11, 6, 'lutff_0/in_3')
// (11, 6, 'sp4_r_v_b_39')
// (11, 7, 'sp12_h_r_23')
// (11, 7, 'sp4_h_r_39')
// (11, 7, 'sp4_r_v_b_26')
// (11, 8, 'local_g2_7')
// (11, 8, 'local_g3_5')
// (11, 8, 'lutff_0/in_3')
// (11, 8, 'lutff_1/in_3')
// (11, 8, 'sp4_r_v_b_15')
// (11, 8, 'sp4_r_v_b_45')
// (11, 9, 'local_g0_3')
// (11, 9, 'lutff_0/in_3')
// (11, 9, 'sp4_r_v_b_2')
// (11, 9, 'sp4_r_v_b_32')
// (11, 10, 'local_g3_5')
// (11, 10, 'lutff_1/in_3')
// (11, 10, 'sp4_r_v_b_21')
// (11, 10, 'sp4_r_v_b_43')
// (11, 11, 'local_g1_6')
// (11, 11, 'lutff_2/in_3')
// (11, 11, 'sp4_r_v_b_30')
// (11, 11, 'sp4_r_v_b_8')
// (11, 12, 'sp4_r_v_b_19')
// (11, 13, 'sp4_r_v_b_6')
// (11, 16, 'neigh_op_tnr_2')
// (11, 16, 'neigh_op_tnr_6')
// (12, 5, 'sp4_v_t_39')
// (12, 6, 'sp4_v_b_39')
// (12, 7, 'sp12_h_l_23')
// (12, 7, 'sp12_v_t_23')
// (12, 7, 'sp4_h_l_39')
// (12, 7, 'sp4_v_b_26')
// (12, 7, 'sp4_v_t_45')
// (12, 8, 'sp12_v_b_23')
// (12, 8, 'sp4_v_b_15')
// (12, 8, 'sp4_v_b_45')
// (12, 9, 'sp12_v_b_20')
// (12, 9, 'sp4_v_b_2')
// (12, 9, 'sp4_v_b_32')
// (12, 9, 'sp4_v_t_43')
// (12, 10, 'sp12_v_b_19')
// (12, 10, 'sp4_v_b_21')
// (12, 10, 'sp4_v_b_43')
// (12, 11, 'sp12_v_b_16')
// (12, 11, 'sp4_v_b_30')
// (12, 11, 'sp4_v_b_8')
// (12, 12, 'sp12_v_b_15')
// (12, 12, 'sp4_v_b_19')
// (12, 13, 'sp12_v_b_12')
// (12, 13, 'sp4_v_b_6')
// (12, 14, 'sp12_v_b_11')
// (12, 15, 'sp12_v_b_8')
// (12, 16, 'neigh_op_top_2')
// (12, 16, 'neigh_op_top_6')
// (12, 16, 'sp12_v_b_7')
// (12, 17, 'io_1/D_IN_0')
// (12, 17, 'io_1/PAD')
// (12, 17, 'span12_vert_4')

wire n27;
// (0, 7, 'span12_horz_4')
// (1, 7, 'sp12_h_r_7')
// (2, 7, 'sp12_h_r_8')
// (3, 7, 'sp12_h_r_11')
// (4, 7, 'sp12_h_r_12')
// (5, 6, 'neigh_op_tnr_4')
// (5, 7, 'neigh_op_rgt_4')
// (5, 7, 'sp12_h_r_15')
// (5, 8, 'neigh_op_bnr_4')
// (6, 6, 'neigh_op_top_4')
// (6, 7, 'lutff_4/out')
// (6, 7, 'sp12_h_r_16')
// (6, 8, 'neigh_op_bot_4')
// (7, 6, 'neigh_op_tnl_4')
// (7, 7, 'local_g0_4')
// (7, 7, 'lutff_0/in_0')
// (7, 7, 'lutff_1/in_3')
// (7, 7, 'neigh_op_lft_4')
// (7, 7, 'sp12_h_r_19')
// (7, 8, 'neigh_op_bnl_4')
// (8, 7, 'local_g0_4')
// (8, 7, 'local_g1_4')
// (8, 7, 'lutff_0/in_1')
// (8, 7, 'lutff_3/in_3')
// (8, 7, 'sp12_h_r_20')
// (9, 7, 'sp12_h_r_23')
// (10, 7, 'sp12_h_l_23')

wire n28;
// (0, 7, 'span12_horz_6')
// (1, 7, 'sp12_h_r_9')
// (2, 7, 'sp12_h_r_10')
// (3, 7, 'sp12_h_r_13')
// (4, 7, 'local_g0_6')
// (4, 7, 'lutff_0/in_2')
// (4, 7, 'sp12_h_r_14')
// (5, 7, 'sp12_h_r_17')
// (6, 7, 'sp12_h_r_18')
// (6, 8, 'sp4_r_v_b_47')
// (6, 9, 'sp4_r_v_b_34')
// (6, 10, 'sp4_r_v_b_23')
// (6, 11, 'sp4_r_v_b_10')
// (7, 6, 'neigh_op_tnr_7')
// (7, 7, 'neigh_op_rgt_7')
// (7, 7, 'sp12_h_r_21')
// (7, 7, 'sp4_h_r_10')
// (7, 7, 'sp4_r_v_b_46')
// (7, 7, 'sp4_v_t_47')
// (7, 8, 'neigh_op_bnr_7')
// (7, 8, 'sp4_r_v_b_35')
// (7, 8, 'sp4_v_b_47')
// (7, 9, 'sp4_r_v_b_22')
// (7, 9, 'sp4_v_b_34')
// (7, 10, 'sp4_r_v_b_11')
// (7, 10, 'sp4_v_b_23')
// (7, 11, 'local_g0_2')
// (7, 11, 'lutff_7/in_3')
// (7, 11, 'sp4_v_b_10')
// (8, 6, 'neigh_op_top_7')
// (8, 6, 'sp4_v_t_46')
// (8, 7, 'lutff_7/out')
// (8, 7, 'sp12_h_r_22')
// (8, 7, 'sp4_h_r_23')
// (8, 7, 'sp4_v_b_46')
// (8, 8, 'local_g0_7')
// (8, 8, 'lutff_0/in_3')
// (8, 8, 'lutff_2/in_3')
// (8, 8, 'neigh_op_bot_7')
// (8, 8, 'sp4_v_b_35')
// (8, 9, 'sp4_v_b_22')
// (8, 10, 'local_g0_3')
// (8, 10, 'local_g1_3')
// (8, 10, 'lutff_0/in_3')
// (8, 10, 'lutff_1/in_3')
// (8, 10, 'lutff_2/in_3')
// (8, 10, 'lutff_7/in_3')
// (8, 10, 'sp4_v_b_11')
// (9, 6, 'neigh_op_tnl_7')
// (9, 7, 'neigh_op_lft_7')
// (9, 7, 'sp12_h_l_22')
// (9, 7, 'sp4_h_r_34')
// (9, 8, 'neigh_op_bnl_7')
// (10, 7, 'sp4_h_r_47')
// (11, 7, 'sp4_h_l_47')

reg n29 = 0;
// (0, 8, 'span12_horz_1')
// (1, 8, 'sp12_h_r_2')
// (2, 8, 'sp12_h_r_5')
// (3, 8, 'sp12_h_r_6')
// (4, 8, 'sp12_h_r_9')
// (5, 8, 'sp12_h_r_10')
// (6, 8, 'sp12_h_r_13')
// (7, 8, 'sp12_h_r_14')
// (8, 7, 'neigh_op_tnr_5')
// (8, 8, 'neigh_op_rgt_5')
// (8, 8, 'sp12_h_r_17')
// (8, 9, 'neigh_op_bnr_5')
// (9, 7, 'neigh_op_top_5')
// (9, 8, 'lutff_5/out')
// (9, 8, 'sp12_h_r_18')
// (9, 9, 'neigh_op_bot_5')
// (10, 7, 'neigh_op_tnl_5')
// (10, 8, 'neigh_op_lft_5')
// (10, 8, 'sp12_h_r_21')
// (10, 9, 'neigh_op_bnl_5')
// (11, 8, 'local_g0_6')
// (11, 8, 'lutff_0/in_2')
// (11, 8, 'sp12_h_r_22')
// (12, 8, 'sp12_h_l_22')

wire n30;
// (0, 8, 'span12_horz_3')
// (1, 8, 'sp12_h_r_4')
// (2, 8, 'sp12_h_r_7')
// (3, 8, 'sp12_h_r_8')
// (4, 8, 'sp12_h_r_11')
// (5, 8, 'sp12_h_r_12')
// (6, 7, 'neigh_op_tnr_4')
// (6, 8, 'neigh_op_rgt_4')
// (6, 8, 'sp12_h_r_15')
// (6, 9, 'neigh_op_bnr_4')
// (7, 7, 'neigh_op_top_4')
// (7, 8, 'lutff_4/out')
// (7, 8, 'sp12_h_r_16')
// (7, 8, 'sp4_h_r_8')
// (7, 9, 'neigh_op_bot_4')
// (8, 7, 'neigh_op_tnl_4')
// (8, 8, 'local_g0_3')
// (8, 8, 'local_g1_5')
// (8, 8, 'lutff_4/in_3')
// (8, 8, 'lutff_6/in_3')
// (8, 8, 'lutff_7/in_3')
// (8, 8, 'neigh_op_lft_4')
// (8, 8, 'sp12_h_r_19')
// (8, 8, 'sp4_h_r_21')
// (8, 9, 'neigh_op_bnl_4')
// (9, 8, 'sp12_h_r_20')
// (9, 8, 'sp4_h_r_32')
// (10, 8, 'sp12_h_r_23')
// (10, 8, 'sp4_h_r_45')
// (11, 8, 'sp12_h_l_23')
// (11, 8, 'sp4_h_l_45')

reg n31 = 0;
// (0, 8, 'span12_horz_6')
// (1, 8, 'sp12_h_r_9')
// (2, 8, 'sp12_h_r_10')
// (3, 7, 'neigh_op_tnr_3')
// (3, 8, 'neigh_op_rgt_3')
// (3, 8, 'sp12_h_r_13')
// (3, 9, 'neigh_op_bnr_3')
// (4, 6, 'sp4_r_v_b_47')
// (4, 7, 'neigh_op_top_3')
// (4, 7, 'sp4_r_v_b_34')
// (4, 8, 'lutff_3/out')
// (4, 8, 'sp12_h_r_14')
// (4, 8, 'sp4_r_v_b_23')
// (4, 8, 'sp4_r_v_b_39')
// (4, 9, 'neigh_op_bot_3')
// (4, 9, 'sp4_r_v_b_10')
// (4, 9, 'sp4_r_v_b_26')
// (4, 10, 'sp4_r_v_b_15')
// (4, 11, 'sp4_r_v_b_2')
// (5, 5, 'sp4_v_t_47')
// (5, 6, 'sp4_v_b_47')
// (5, 7, 'neigh_op_tnl_3')
// (5, 7, 'sp4_v_b_34')
// (5, 7, 'sp4_v_t_39')
// (5, 8, 'neigh_op_lft_3')
// (5, 8, 'sp12_h_r_17')
// (5, 8, 'sp4_v_b_23')
// (5, 8, 'sp4_v_b_39')
// (5, 9, 'neigh_op_bnl_3')
// (5, 9, 'sp4_h_r_10')
// (5, 9, 'sp4_v_b_10')
// (5, 9, 'sp4_v_b_26')
// (5, 10, 'sp4_v_b_15')
// (5, 11, 'sp4_h_r_11')
// (5, 11, 'sp4_h_r_8')
// (5, 11, 'sp4_v_b_2')
// (6, 8, 'sp12_h_r_18')
// (6, 9, 'sp4_h_r_23')
// (6, 11, 'sp4_h_r_21')
// (6, 11, 'sp4_h_r_22')
// (7, 8, 'sp12_h_r_21')
// (7, 8, 'sp4_h_r_10')
// (7, 9, 'sp4_h_r_34')
// (7, 11, 'local_g2_0')
// (7, 11, 'local_g2_3')
// (7, 11, 'lutff_4/in_2')
// (7, 11, 'lutff_7/in_2')
// (7, 11, 'sp4_h_r_32')
// (7, 11, 'sp4_h_r_35')
// (8, 8, 'sp12_h_r_22')
// (8, 8, 'sp4_h_r_23')
// (8, 8, 'sp4_r_v_b_45')
// (8, 8, 'sp4_r_v_b_46')
// (8, 9, 'local_g0_3')
// (8, 9, 'local_g2_0')
// (8, 9, 'lutff_2/in_0')
// (8, 9, 'lutff_3/in_2')
// (8, 9, 'lutff_4/in_2')
// (8, 9, 'lutff_6/in_1')
// (8, 9, 'sp4_h_r_47')
// (8, 9, 'sp4_r_v_b_32')
// (8, 9, 'sp4_r_v_b_35')
// (8, 10, 'local_g3_5')
// (8, 10, 'local_g3_6')
// (8, 10, 'lutff_0/in_2')
// (8, 10, 'lutff_1/in_0')
// (8, 10, 'lutff_2/in_2')
// (8, 10, 'lutff_6/in_2')
// (8, 10, 'lutff_7/in_0')
// (8, 10, 'sp4_r_v_b_21')
// (8, 10, 'sp4_r_v_b_22')
// (8, 11, 'local_g3_5')
// (8, 11, 'lutff_2/in_2')
// (8, 11, 'sp4_h_r_45')
// (8, 11, 'sp4_h_r_46')
// (8, 11, 'sp4_r_v_b_11')
// (8, 11, 'sp4_r_v_b_8')
// (8, 12, 'sp4_r_v_b_46')
// (8, 13, 'local_g0_0')
// (8, 13, 'local_g2_3')
// (8, 13, 'lutff_1/in_2')
// (8, 13, 'lutff_3/in_2')
// (8, 13, 'lutff_4/in_0')
// (8, 13, 'lutff_6/in_2')
// (8, 13, 'sp4_r_v_b_35')
// (8, 14, 'sp4_r_v_b_22')
// (8, 15, 'sp4_r_v_b_11')
// (9, 7, 'sp4_v_t_45')
// (9, 7, 'sp4_v_t_46')
// (9, 8, 'sp12_h_l_22')
// (9, 8, 'sp4_h_r_34')
// (9, 8, 'sp4_v_b_45')
// (9, 8, 'sp4_v_b_46')
// (9, 9, 'local_g2_0')
// (9, 9, 'local_g3_0')
// (9, 9, 'lutff_2/in_0')
// (9, 9, 'lutff_4/in_2')
// (9, 9, 'lutff_5/in_2')
// (9, 9, 'lutff_7/in_2')
// (9, 9, 'sp4_h_l_47')
// (9, 9, 'sp4_h_r_1')
// (9, 9, 'sp4_v_b_32')
// (9, 9, 'sp4_v_b_35')
// (9, 10, 'sp4_v_b_21')
// (9, 10, 'sp4_v_b_22')
// (9, 11, 'sp4_h_l_45')
// (9, 11, 'sp4_h_l_46')
// (9, 11, 'sp4_v_b_11')
// (9, 11, 'sp4_v_b_8')
// (9, 11, 'sp4_v_t_46')
// (9, 12, 'local_g2_6')
// (9, 12, 'local_g3_6')
// (9, 12, 'lutff_1/in_2')
// (9, 12, 'lutff_6/in_2')
// (9, 12, 'lutff_7/in_2')
// (9, 12, 'sp4_v_b_46')
// (9, 13, 'sp4_v_b_35')
// (9, 14, 'sp4_v_b_22')
// (9, 15, 'sp4_v_b_11')
// (10, 8, 'sp4_h_r_47')
// (10, 9, 'sp4_h_r_12')
// (10, 9, 'sp4_r_v_b_38')
// (10, 9, 'sp4_r_v_b_47')
// (10, 10, 'sp4_r_v_b_27')
// (10, 10, 'sp4_r_v_b_34')
// (10, 11, 'sp4_r_v_b_14')
// (10, 11, 'sp4_r_v_b_23')
// (10, 12, 'sp4_r_v_b_10')
// (10, 12, 'sp4_r_v_b_3')
// (11, 8, 'sp4_h_l_47')
// (11, 8, 'sp4_v_t_38')
// (11, 8, 'sp4_v_t_47')
// (11, 9, 'local_g2_1')
// (11, 9, 'local_g3_1')
// (11, 9, 'lutff_1/in_2')
// (11, 9, 'lutff_4/in_0')
// (11, 9, 'lutff_5/in_2')
// (11, 9, 'lutff_6/in_2')
// (11, 9, 'sp4_h_r_25')
// (11, 9, 'sp4_v_b_38')
// (11, 9, 'sp4_v_b_47')
// (11, 10, 'sp4_v_b_27')
// (11, 10, 'sp4_v_b_34')
// (11, 11, 'sp4_v_b_14')
// (11, 11, 'sp4_v_b_23')
// (11, 12, 'local_g0_2')
// (11, 12, 'local_g0_3')
// (11, 12, 'lutff_0/in_1')
// (11, 12, 'lutff_1/in_2')
// (11, 12, 'lutff_3/in_2')
// (11, 12, 'lutff_6/in_2')
// (11, 12, 'lutff_7/in_0')
// (11, 12, 'sp4_v_b_10')
// (11, 12, 'sp4_v_b_3')
// (12, 9, 'sp4_h_r_36')
// (13, 9, 'span4_horz_36')

reg n32 = 0;
// (0, 9, 'span12_horz_1')
// (1, 9, 'sp12_h_r_2')
// (2, 9, 'sp12_h_r_5')
// (3, 9, 'sp12_h_r_6')
// (4, 9, 'sp12_h_r_9')
// (5, 9, 'sp12_h_r_10')
// (6, 8, 'neigh_op_tnr_3')
// (6, 9, 'neigh_op_rgt_3')
// (6, 9, 'sp12_h_r_13')
// (6, 10, 'neigh_op_bnr_3')
// (7, 5, 'sp4_r_v_b_40')
// (7, 6, 'local_g1_5')
// (7, 6, 'lutff_1/in_3')
// (7, 6, 'sp4_r_v_b_29')
// (7, 7, 'sp4_r_v_b_16')
// (7, 8, 'neigh_op_top_3')
// (7, 8, 'sp4_r_v_b_5')
// (7, 9, 'lutff_3/out')
// (7, 9, 'sp12_h_r_14')
// (7, 9, 'sp4_r_v_b_39')
// (7, 10, 'neigh_op_bot_3')
// (7, 10, 'sp4_r_v_b_26')
// (7, 11, 'sp4_r_v_b_15')
// (7, 12, 'sp4_r_v_b_2')
// (8, 4, 'sp4_v_t_40')
// (8, 5, 'sp4_v_b_40')
// (8, 6, 'sp4_v_b_29')
// (8, 7, 'sp4_v_b_16')
// (8, 8, 'neigh_op_tnl_3')
// (8, 8, 'sp4_v_b_5')
// (8, 8, 'sp4_v_t_39')
// (8, 9, 'neigh_op_lft_3')
// (8, 9, 'sp12_h_r_17')
// (8, 9, 'sp4_v_b_39')
// (8, 10, 'neigh_op_bnl_3')
// (8, 10, 'sp4_v_b_26')
// (8, 11, 'sp4_v_b_15')
// (8, 12, 'sp4_v_b_2')
// (9, 9, 'sp12_h_r_18')
// (10, 9, 'sp12_h_r_21')
// (11, 9, 'local_g1_6')
// (11, 9, 'lutff_0/in_1')
// (11, 9, 'sp12_h_r_22')
// (12, 9, 'sp12_h_l_22')

reg n33 = 0;
// (0, 9, 'span12_horz_10')
// (1, 8, 'neigh_op_tnr_3')
// (1, 9, 'neigh_op_rgt_3')
// (1, 9, 'sp12_h_r_13')
// (1, 10, 'neigh_op_bnr_3')
// (2, 8, 'neigh_op_top_3')
// (2, 9, 'lutff_3/out')
// (2, 9, 'sp12_h_r_14')
// (2, 10, 'neigh_op_bot_3')
// (3, 8, 'neigh_op_tnl_3')
// (3, 9, 'neigh_op_lft_3')
// (3, 9, 'sp12_h_r_17')
// (3, 10, 'neigh_op_bnl_3')
// (4, 9, 'sp12_h_r_18')
// (5, 9, 'local_g1_5')
// (5, 9, 'lutff_4/in_0')
// (5, 9, 'sp12_h_r_21')
// (6, 9, 'sp12_h_r_22')
// (7, 9, 'sp12_h_l_22')

reg n34 = 0;
// (0, 9, 'span12_horz_2')
// (1, 9, 'sp12_h_r_5')
// (2, 9, 'local_g0_6')
// (2, 9, 'lutff_2/in_0')
// (2, 9, 'sp12_h_r_6')
// (3, 8, 'neigh_op_tnr_1')
// (3, 9, 'neigh_op_rgt_1')
// (3, 9, 'sp12_h_r_9')
// (3, 10, 'neigh_op_bnr_1')
// (4, 8, 'neigh_op_top_1')
// (4, 9, 'lutff_1/out')
// (4, 9, 'sp12_h_r_10')
// (4, 10, 'neigh_op_bot_1')
// (5, 8, 'neigh_op_tnl_1')
// (5, 9, 'neigh_op_lft_1')
// (5, 9, 'sp12_h_r_13')
// (5, 10, 'neigh_op_bnl_1')
// (6, 9, 'sp12_h_r_14')
// (7, 9, 'sp12_h_r_17')
// (8, 9, 'sp12_h_r_18')
// (9, 9, 'sp12_h_r_21')
// (10, 9, 'sp12_h_r_22')
// (11, 9, 'sp12_h_l_22')

reg n35 = 0;
// (0, 9, 'span12_horz_4')
// (1, 9, 'sp12_h_r_7')
// (2, 9, 'sp12_h_r_8')
// (3, 8, 'neigh_op_tnr_2')
// (3, 9, 'neigh_op_rgt_2')
// (3, 9, 'sp12_h_r_11')
// (3, 10, 'neigh_op_bnr_2')
// (4, 8, 'neigh_op_top_2')
// (4, 9, 'lutff_2/out')
// (4, 9, 'sp12_h_r_12')
// (4, 10, 'neigh_op_bot_2')
// (5, 8, 'neigh_op_tnl_2')
// (5, 9, 'neigh_op_lft_2')
// (5, 9, 'sp12_h_r_15')
// (5, 10, 'neigh_op_bnl_2')
// (6, 9, 'sp12_h_r_16')
// (7, 9, 'local_g0_3')
// (7, 9, 'lutff_2/in_3')
// (7, 9, 'sp12_h_r_19')
// (8, 9, 'sp12_h_r_20')
// (9, 9, 'sp12_h_r_23')
// (10, 9, 'sp12_h_l_23')

reg n36 = 0;
// (0, 9, 'span12_horz_6')
// (1, 9, 'sp12_h_r_9')
// (2, 9, 'local_g0_2')
// (2, 9, 'lutff_0/in_0')
// (2, 9, 'sp12_h_r_10')
// (3, 8, 'neigh_op_tnr_3')
// (3, 9, 'neigh_op_rgt_3')
// (3, 9, 'sp12_h_r_13')
// (3, 10, 'neigh_op_bnr_3')
// (4, 8, 'neigh_op_top_3')
// (4, 9, 'lutff_3/out')
// (4, 9, 'sp12_h_r_14')
// (4, 10, 'neigh_op_bot_3')
// (5, 8, 'neigh_op_tnl_3')
// (5, 9, 'neigh_op_lft_3')
// (5, 9, 'sp12_h_r_17')
// (5, 10, 'neigh_op_bnl_3')
// (6, 9, 'sp12_h_r_18')
// (7, 9, 'sp12_h_r_21')
// (8, 9, 'sp12_h_r_22')
// (9, 9, 'sp12_h_l_22')

reg n37 = 0;
// (0, 10, 'span12_horz_5')
// (1, 10, 'sp12_h_r_6')
// (2, 10, 'sp12_h_r_9')
// (3, 10, 'sp12_h_r_10')
// (4, 9, 'neigh_op_tnr_3')
// (4, 10, 'neigh_op_rgt_3')
// (4, 10, 'sp12_h_r_13')
// (4, 11, 'neigh_op_bnr_3')
// (5, 3, 'sp4_r_v_b_42')
// (5, 4, 'sp4_r_v_b_31')
// (5, 5, 'sp4_r_v_b_18')
// (5, 6, 'sp4_r_v_b_7')
// (5, 7, 'sp4_r_v_b_42')
// (5, 8, 'sp4_r_v_b_31')
// (5, 9, 'neigh_op_top_3')
// (5, 9, 'sp4_r_v_b_18')
// (5, 10, 'lutff_3/out')
// (5, 10, 'sp12_h_r_14')
// (5, 10, 'sp4_r_v_b_7')
// (5, 11, 'neigh_op_bot_3')
// (6, 2, 'sp4_v_t_42')
// (6, 3, 'sp4_v_b_42')
// (6, 4, 'sp4_v_b_31')
// (6, 5, 'sp4_v_b_18')
// (6, 6, 'sp4_h_r_1')
// (6, 6, 'sp4_v_b_7')
// (6, 6, 'sp4_v_t_42')
// (6, 7, 'sp4_v_b_42')
// (6, 8, 'sp4_v_b_31')
// (6, 9, 'neigh_op_tnl_3')
// (6, 9, 'sp4_v_b_18')
// (6, 10, 'neigh_op_lft_3')
// (6, 10, 'sp12_h_r_17')
// (6, 10, 'sp4_v_b_7')
// (6, 11, 'neigh_op_bnl_3')
// (7, 6, 'local_g1_4')
// (7, 6, 'lutff_0/in_3')
// (7, 6, 'sp4_h_r_12')
// (7, 10, 'sp12_h_r_18')
// (8, 6, 'sp4_h_r_25')
// (8, 10, 'sp12_h_r_21')
// (9, 6, 'sp4_h_r_36')
// (9, 10, 'sp12_h_r_22')
// (10, 6, 'sp4_h_l_36')
// (10, 10, 'sp12_h_l_22')
// (10, 10, 'sp12_h_r_1')
// (11, 10, 'local_g0_2')
// (11, 10, 'lutff_1/in_1')
// (11, 10, 'sp12_h_r_2')
// (12, 10, 'sp12_h_r_5')
// (13, 10, 'span12_horz_5')

wire n38;
// (0, 10, 'span12_horz_6')
// (1, 10, 'sp12_h_r_9')
// (2, 10, 'sp12_h_r_10')
// (3, 10, 'sp12_h_r_13')
// (4, 10, 'sp12_h_r_14')
// (5, 10, 'local_g0_1')
// (5, 10, 'local_g1_1')
// (5, 10, 'lutff_2/in_1')
// (5, 10, 'lutff_7/in_1')
// (5, 10, 'sp12_h_r_17')
// (6, 10, 'sp12_h_r_18')
// (7, 10, 'sp12_h_r_21')
// (8, 8, 'neigh_op_tnr_1')
// (8, 9, 'neigh_op_rgt_1')
// (8, 10, 'neigh_op_bnr_1')
// (8, 10, 'sp12_h_r_22')
// (9, 0, 'span12_vert_18')
// (9, 1, 'sp12_v_b_18')
// (9, 2, 'sp12_v_b_17')
// (9, 3, 'sp12_v_b_14')
// (9, 4, 'sp12_v_b_13')
// (9, 5, 'sp12_v_b_10')
// (9, 6, 'sp12_v_b_9')
// (9, 7, 'sp12_v_b_6')
// (9, 8, 'neigh_op_top_1')
// (9, 8, 'sp12_v_b_5')
// (9, 9, 'lutff_1/out')
// (9, 9, 'sp12_v_b_2')
// (9, 10, 'neigh_op_bot_1')
// (9, 10, 'sp12_h_l_22')
// (9, 10, 'sp12_v_b_1')
// (10, 8, 'neigh_op_tnl_1')
// (10, 9, 'neigh_op_lft_1')
// (10, 10, 'neigh_op_bnl_1')

reg n39 = 0;
// (0, 10, 'span12_horz_7')
// (1, 10, 'sp12_h_r_8')
// (2, 10, 'sp12_h_r_11')
// (3, 10, 'sp12_h_r_12')
// (4, 10, 'sp12_h_r_15')
// (5, 10, 'sp12_h_r_16')
// (6, 9, 'neigh_op_tnr_6')
// (6, 10, 'neigh_op_rgt_6')
// (6, 10, 'sp12_h_r_19')
// (6, 11, 'neigh_op_bnr_6')
// (7, 9, 'neigh_op_top_6')
// (7, 10, 'lutff_6/out')
// (7, 10, 'sp12_h_r_20')
// (7, 11, 'neigh_op_bot_6')
// (8, 9, 'neigh_op_tnl_6')
// (8, 10, 'neigh_op_lft_6')
// (8, 10, 'sp12_h_r_23')
// (8, 11, 'neigh_op_bnl_6')
// (9, 0, 'span12_vert_19')
// (9, 1, 'sp12_v_b_19')
// (9, 2, 'sp12_v_b_16')
// (9, 3, 'sp12_v_b_15')
// (9, 4, 'sp12_v_b_12')
// (9, 5, 'local_g3_3')
// (9, 5, 'lutff_4/in_0')
// (9, 5, 'sp12_v_b_11')
// (9, 6, 'sp12_v_b_8')
// (9, 7, 'sp12_v_b_7')
// (9, 8, 'sp12_v_b_4')
// (9, 9, 'sp12_v_b_3')
// (9, 10, 'sp12_h_l_23')
// (9, 10, 'sp12_v_b_0')

reg n40 = 0;
// (0, 10, 'span4_horz_8')
// (1, 9, 'neigh_op_tnr_0')
// (1, 10, 'neigh_op_rgt_0')
// (1, 10, 'sp4_h_r_21')
// (1, 11, 'neigh_op_bnr_0')
// (2, 9, 'neigh_op_top_0')
// (2, 10, 'lutff_0/out')
// (2, 10, 'sp4_h_r_32')
// (2, 11, 'neigh_op_bot_0')
// (3, 7, 'sp4_r_v_b_39')
// (3, 8, 'sp4_r_v_b_26')
// (3, 9, 'neigh_op_tnl_0')
// (3, 9, 'sp4_r_v_b_15')
// (3, 10, 'neigh_op_lft_0')
// (3, 10, 'sp4_h_r_45')
// (3, 10, 'sp4_r_v_b_2')
// (3, 11, 'neigh_op_bnl_0')
// (4, 6, 'sp4_v_t_39')
// (4, 7, 'sp4_v_b_39')
// (4, 8, 'sp4_v_b_26')
// (4, 9, 'local_g1_7')
// (4, 9, 'lutff_2/in_0')
// (4, 9, 'sp4_v_b_15')
// (4, 10, 'sp4_h_l_45')
// (4, 10, 'sp4_v_b_2')

reg n41 = 0;
// (0, 12, 'span12_horz_1')
// (1, 12, 'sp12_h_r_2')
// (2, 12, 'sp12_h_r_5')
// (3, 12, 'sp12_h_r_6')
// (4, 12, 'sp12_h_r_9')
// (5, 12, 'sp12_h_r_10')
// (6, 12, 'sp12_h_r_13')
// (7, 12, 'sp12_h_r_14')
// (8, 12, 'sp12_h_r_17')
// (9, 12, 'local_g1_2')
// (9, 12, 'lutff_3/in_2')
// (9, 12, 'sp12_h_r_18')
// (10, 11, 'neigh_op_tnr_7')
// (10, 12, 'neigh_op_rgt_7')
// (10, 12, 'sp12_h_r_21')
// (10, 13, 'neigh_op_bnr_7')
// (11, 11, 'neigh_op_top_7')
// (11, 12, 'local_g0_7')
// (11, 12, 'lutff_6/in_1')
// (11, 12, 'lutff_7/out')
// (11, 12, 'sp12_h_r_22')
// (11, 13, 'neigh_op_bot_7')
// (12, 11, 'neigh_op_tnl_7')
// (12, 12, 'neigh_op_lft_7')
// (12, 12, 'sp12_h_l_22')
// (12, 13, 'neigh_op_bnl_7')

reg n42 = 0;
// (0, 12, 'span12_horz_8')
// (1, 12, 'sp12_h_r_11')
// (2, 12, 'sp12_h_r_12')
// (3, 12, 'sp12_h_r_15')
// (4, 12, 'sp12_h_r_16')
// (5, 11, 'neigh_op_tnr_6')
// (5, 12, 'neigh_op_rgt_6')
// (5, 12, 'sp12_h_r_19')
// (5, 13, 'neigh_op_bnr_6')
// (6, 11, 'neigh_op_top_6')
// (6, 12, 'lutff_6/out')
// (6, 12, 'sp12_h_r_20')
// (6, 13, 'neigh_op_bot_6')
// (7, 11, 'neigh_op_tnl_6')
// (7, 12, 'local_g0_7')
// (7, 12, 'lutff_3/in_0')
// (7, 12, 'neigh_op_lft_6')
// (7, 12, 'sp12_h_r_23')
// (7, 13, 'neigh_op_bnl_6')
// (8, 12, 'sp12_h_l_23')

reg n43 = 0;
// (0, 13, 'span12_horz_1')
// (1, 13, 'sp12_h_r_2')
// (2, 13, 'sp12_h_r_5')
// (3, 13, 'sp12_h_r_6')
// (4, 13, 'sp12_h_r_9')
// (5, 12, 'sp4_r_v_b_38')
// (5, 13, 'sp12_h_r_10')
// (5, 13, 'sp4_r_v_b_27')
// (5, 14, 'sp4_r_v_b_14')
// (5, 15, 'sp4_r_v_b_3')
// (6, 11, 'local_g1_1')
// (6, 11, 'lutff_4/in_0')
// (6, 11, 'sp4_h_r_9')
// (6, 11, 'sp4_v_t_38')
// (6, 12, 'local_g2_6')
// (6, 12, 'local_g3_6')
// (6, 12, 'lutff_3/in_0')
// (6, 12, 'lutff_6/in_0')
// (6, 12, 'sp4_v_b_38')
// (6, 13, 'sp12_h_r_13')
// (6, 13, 'sp4_v_b_27')
// (6, 14, 'sp4_v_b_14')
// (6, 15, 'sp4_v_b_3')
// (7, 11, 'sp4_h_r_20')
// (7, 13, 'local_g1_6')
// (7, 13, 'lutff_3/in_0')
// (7, 13, 'sp12_h_r_14')
// (8, 11, 'sp4_h_r_33')
// (8, 12, 'neigh_op_tnr_5')
// (8, 13, 'neigh_op_rgt_5')
// (8, 13, 'sp12_h_r_17')
// (8, 14, 'neigh_op_bnr_5')
// (9, 11, 'sp4_h_r_44')
// (9, 12, 'neigh_op_top_5')
// (9, 12, 'sp4_r_v_b_38')
// (9, 13, 'lutff_5/out')
// (9, 13, 'sp12_h_r_18')
// (9, 13, 'sp4_r_v_b_27')
// (9, 14, 'neigh_op_bot_5')
// (9, 14, 'sp4_r_v_b_14')
// (9, 15, 'sp4_r_v_b_3')
// (10, 11, 'sp4_h_l_44')
// (10, 11, 'sp4_v_t_38')
// (10, 12, 'neigh_op_tnl_5')
// (10, 12, 'sp4_v_b_38')
// (10, 13, 'neigh_op_lft_5')
// (10, 13, 'sp12_h_r_21')
// (10, 13, 'sp4_v_b_27')
// (10, 14, 'neigh_op_bnl_5')
// (10, 14, 'sp4_v_b_14')
// (10, 15, 'sp4_v_b_3')
// (11, 13, 'sp12_h_r_22')
// (12, 13, 'sp12_h_l_22')

reg d_vld = 0;
// (0, 14, 'io_0/D_OUT_0')
// (0, 14, 'io_0/PAD')
// (0, 14, 'local_g0_0')
// (0, 14, 'span4_horz_24')
// (1, 7, 'neigh_op_tnr_3')
// (1, 8, 'neigh_op_rgt_3')
// (1, 9, 'neigh_op_bnr_3')
// (1, 11, 'sp4_r_v_b_42')
// (1, 12, 'sp4_r_v_b_31')
// (1, 13, 'sp4_r_v_b_18')
// (1, 14, 'sp4_h_r_37')
// (1, 14, 'sp4_r_v_b_7')
// (2, 7, 'neigh_op_top_3')
// (2, 7, 'sp12_v_t_22')
// (2, 8, 'lutff_3/out')
// (2, 8, 'sp12_v_b_22')
// (2, 9, 'neigh_op_bot_3')
// (2, 9, 'sp12_v_b_21')
// (2, 10, 'sp12_v_b_18')
// (2, 10, 'sp4_v_t_42')
// (2, 11, 'sp12_v_b_17')
// (2, 11, 'sp4_v_b_42')
// (2, 12, 'sp12_v_b_14')
// (2, 12, 'sp4_v_b_31')
// (2, 13, 'sp12_v_b_13')
// (2, 13, 'sp4_v_b_18')
// (2, 14, 'sp12_v_b_10')
// (2, 14, 'sp4_h_l_37')
// (2, 14, 'sp4_v_b_7')
// (2, 15, 'sp12_v_b_9')
// (2, 16, 'sp12_v_b_6')
// (2, 17, 'span12_vert_5')
// (3, 7, 'neigh_op_tnl_3')
// (3, 8, 'neigh_op_lft_3')
// (3, 9, 'neigh_op_bnl_3')

reg n45 = 0;
// (0, 14, 'span12_horz_10')
// (1, 13, 'neigh_op_tnr_3')
// (1, 14, 'neigh_op_rgt_3')
// (1, 14, 'sp12_h_r_13')
// (1, 15, 'neigh_op_bnr_3')
// (2, 13, 'neigh_op_top_3')
// (2, 14, 'lutff_3/out')
// (2, 14, 'sp12_h_r_14')
// (2, 15, 'neigh_op_bot_3')
// (3, 13, 'neigh_op_tnl_3')
// (3, 14, 'neigh_op_lft_3')
// (3, 14, 'sp12_h_r_17')
// (3, 15, 'neigh_op_bnl_3')
// (4, 14, 'local_g1_2')
// (4, 14, 'lutff_3/in_0')
// (4, 14, 'sp12_h_r_18')
// (5, 14, 'sp12_h_r_21')
// (6, 14, 'sp12_h_r_22')
// (7, 14, 'sp12_h_l_22')

reg n46 = 0;
// (0, 14, 'span12_horz_6')
// (1, 14, 'sp12_h_r_9')
// (2, 14, 'sp12_h_r_10')
// (3, 13, 'neigh_op_tnr_3')
// (3, 14, 'neigh_op_rgt_3')
// (3, 14, 'sp12_h_r_13')
// (3, 15, 'neigh_op_bnr_3')
// (4, 13, 'neigh_op_top_3')
// (4, 14, 'lutff_3/out')
// (4, 14, 'sp12_h_r_14')
// (4, 15, 'neigh_op_bot_3')
// (5, 13, 'neigh_op_tnl_3')
// (5, 14, 'local_g1_1')
// (5, 14, 'lutff_0/in_0')
// (5, 14, 'neigh_op_lft_3')
// (5, 14, 'sp12_h_r_17')
// (5, 15, 'neigh_op_bnl_3')
// (6, 14, 'sp12_h_r_18')
// (7, 14, 'sp12_h_r_21')
// (8, 14, 'sp12_h_r_22')
// (9, 14, 'sp12_h_l_22')

reg n47 = 0;
// (0, 14, 'span12_horz_7')
// (1, 14, 'sp12_h_r_8')
// (2, 14, 'local_g0_3')
// (2, 14, 'lutff_3/in_0')
// (2, 14, 'sp12_h_r_11')
// (3, 14, 'sp12_h_r_12')
// (4, 13, 'neigh_op_tnr_4')
// (4, 14, 'neigh_op_rgt_4')
// (4, 14, 'sp12_h_r_15')
// (4, 15, 'neigh_op_bnr_4')
// (5, 13, 'neigh_op_top_4')
// (5, 14, 'lutff_4/out')
// (5, 14, 'sp12_h_r_16')
// (5, 15, 'neigh_op_bot_4')
// (6, 13, 'neigh_op_tnl_4')
// (6, 14, 'neigh_op_lft_4')
// (6, 14, 'sp12_h_r_19')
// (6, 15, 'neigh_op_bnl_4')
// (7, 14, 'sp12_h_r_20')
// (8, 14, 'sp12_h_r_23')
// (9, 14, 'sp12_h_l_23')

wire n48;
// (1, 1, 'neigh_op_tnr_1')
// (1, 2, 'neigh_op_rgt_1')
// (1, 3, 'neigh_op_bnr_1')
// (2, 1, 'neigh_op_top_1')
// (2, 1, 'sp4_r_v_b_46')
// (2, 2, 'local_g1_1')
// (2, 2, 'lutff_1/out')
// (2, 2, 'lutff_2/in_2')
// (2, 2, 'sp4_r_v_b_35')
// (2, 3, 'local_g3_6')
// (2, 3, 'lutff_1/in_2')
// (2, 3, 'neigh_op_bot_1')
// (2, 3, 'sp4_r_v_b_22')
// (2, 4, 'sp4_r_v_b_11')
// (3, 0, 'span4_vert_46')
// (3, 1, 'neigh_op_tnl_1')
// (3, 1, 'sp4_v_b_46')
// (3, 2, 'neigh_op_lft_1')
// (3, 2, 'sp4_v_b_35')
// (3, 3, 'neigh_op_bnl_1')
// (3, 3, 'sp4_v_b_22')
// (3, 4, 'sp4_v_b_11')

reg n49 = 0;
// (1, 1, 'neigh_op_tnr_2')
// (1, 2, 'neigh_op_rgt_2')
// (1, 2, 'sp4_h_r_9')
// (1, 2, 'sp4_r_v_b_36')
// (1, 3, 'neigh_op_bnr_2')
// (1, 3, 'sp4_r_v_b_25')
// (1, 4, 'sp4_r_v_b_12')
// (1, 5, 'sp4_r_v_b_1')
// (2, 1, 'neigh_op_top_2')
// (2, 1, 'sp4_v_t_36')
// (2, 2, 'local_g0_2')
// (2, 2, 'lutff_1/in_3')
// (2, 2, 'lutff_2/out')
// (2, 2, 'sp4_h_r_20')
// (2, 2, 'sp4_v_b_36')
// (2, 3, 'neigh_op_bot_2')
// (2, 3, 'sp4_v_b_25')
// (2, 4, 'local_g1_4')
// (2, 4, 'lutff_7/in_2')
// (2, 4, 'sp4_v_b_12')
// (2, 5, 'sp4_h_r_10')
// (2, 5, 'sp4_h_r_7')
// (2, 5, 'sp4_v_b_1')
// (3, 1, 'neigh_op_tnl_2')
// (3, 2, 'neigh_op_lft_2')
// (3, 2, 'sp4_h_r_33')
// (3, 3, 'neigh_op_bnl_2')
// (3, 5, 'sp4_h_r_18')
// (3, 5, 'sp4_h_r_23')
// (4, 2, 'local_g2_4')
// (4, 2, 'lutff_5/in_3')
// (4, 2, 'sp4_h_r_44')
// (4, 3, 'sp4_r_v_b_39')
// (4, 4, 'sp4_r_v_b_26')
// (4, 5, 'sp4_h_r_31')
// (4, 5, 'sp4_h_r_34')
// (4, 5, 'sp4_r_v_b_15')
// (4, 6, 'sp4_r_v_b_2')
// (5, 2, 'sp4_h_l_44')
// (5, 2, 'sp4_h_r_5')
// (5, 2, 'sp4_r_v_b_36')
// (5, 2, 'sp4_r_v_b_41')
// (5, 2, 'sp4_v_t_39')
// (5, 3, 'sp4_r_v_b_25')
// (5, 3, 'sp4_r_v_b_28')
// (5, 3, 'sp4_v_b_39')
// (5, 4, 'local_g2_2')
// (5, 4, 'lutff_0/in_0')
// (5, 4, 'lutff_4/in_0')
// (5, 4, 'sp4_r_v_b_12')
// (5, 4, 'sp4_r_v_b_17')
// (5, 4, 'sp4_v_b_26')
// (5, 5, 'local_g1_7')
// (5, 5, 'local_g3_2')
// (5, 5, 'lutff_0/in_0')
// (5, 5, 'lutff_1/in_0')
// (5, 5, 'lutff_2/in_0')
// (5, 5, 'lutff_4/in_0')
// (5, 5, 'lutff_5/in_0')
// (5, 5, 'sp4_h_r_42')
// (5, 5, 'sp4_h_r_47')
// (5, 5, 'sp4_r_v_b_1')
// (5, 5, 'sp4_r_v_b_4')
// (5, 5, 'sp4_v_b_15')
// (5, 6, 'sp4_v_b_2')
// (6, 1, 'sp4_v_t_36')
// (6, 1, 'sp4_v_t_41')
// (6, 2, 'local_g0_0')
// (6, 2, 'lutff_2/in_2')
// (6, 2, 'sp4_h_r_16')
// (6, 2, 'sp4_v_b_36')
// (6, 2, 'sp4_v_b_41')
// (6, 3, 'local_g3_1')
// (6, 3, 'lutff_2/in_0')
// (6, 3, 'lutff_4/in_0')
// (6, 3, 'sp4_v_b_25')
// (6, 3, 'sp4_v_b_28')
// (6, 4, 'local_g0_1')
// (6, 4, 'lutff_3/in_0')
// (6, 4, 'sp4_v_b_12')
// (6, 4, 'sp4_v_b_17')
// (6, 5, 'local_g0_2')
// (6, 5, 'local_g1_6')
// (6, 5, 'lutff_0/in_0')
// (6, 5, 'lutff_1/in_0')
// (6, 5, 'lutff_2/in_0')
// (6, 5, 'lutff_3/in_1')
// (6, 5, 'lutff_4/in_0')
// (6, 5, 'sp4_h_l_42')
// (6, 5, 'sp4_h_l_47')
// (6, 5, 'sp4_h_r_10')
// (6, 5, 'sp4_h_r_6')
// (6, 5, 'sp4_v_b_1')
// (6, 5, 'sp4_v_b_4')
// (7, 2, 'sp4_h_r_29')
// (7, 5, 'sp4_h_r_19')
// (7, 5, 'sp4_h_r_23')
// (8, 2, 'sp4_h_r_40')
// (8, 5, 'sp4_h_r_30')
// (8, 5, 'sp4_h_r_34')
// (9, 2, 'sp4_h_l_40')
// (9, 5, 'sp4_h_r_43')
// (9, 5, 'sp4_h_r_47')
// (10, 5, 'sp4_h_l_43')
// (10, 5, 'sp4_h_l_47')

wire n50;
// (1, 2, 'neigh_op_tnr_0')
// (1, 3, 'neigh_op_rgt_0')
// (1, 4, 'neigh_op_bnr_0')
// (2, 2, 'local_g0_0')
// (2, 2, 'lutff_2/in_0')
// (2, 2, 'lutff_4/in_0')
// (2, 2, 'neigh_op_top_0')
// (2, 3, 'local_g0_0')
// (2, 3, 'lutff_0/out')
// (2, 3, 'lutff_4/in_2')
// (2, 4, 'neigh_op_bot_0')
// (3, 2, 'neigh_op_tnl_0')
// (3, 3, 'neigh_op_lft_0')
// (3, 4, 'neigh_op_bnl_0')

wire n51;
// (1, 2, 'neigh_op_tnr_1')
// (1, 3, 'local_g2_1')
// (1, 3, 'local_g3_1')
// (1, 3, 'lutff_2/in_0')
// (1, 3, 'lutff_3/in_0')
// (1, 3, 'lutff_4/in_0')
// (1, 3, 'neigh_op_rgt_1')
// (1, 4, 'neigh_op_bnr_1')
// (2, 2, 'neigh_op_top_1')
// (2, 3, 'lutff_1/out')
// (2, 4, 'neigh_op_bot_1')
// (3, 2, 'neigh_op_tnl_1')
// (3, 3, 'neigh_op_lft_1')
// (3, 4, 'neigh_op_bnl_1')

wire n52;
// (1, 2, 'neigh_op_tnr_2')
// (1, 3, 'neigh_op_rgt_2')
// (1, 3, 'sp4_r_v_b_36')
// (1, 4, 'neigh_op_bnr_2')
// (1, 4, 'sp4_r_v_b_25')
// (1, 5, 'sp4_r_v_b_12')
// (1, 6, 'sp4_r_v_b_1')
// (2, 2, 'local_g1_2')
// (2, 2, 'lutff_6/in_1')
// (2, 2, 'neigh_op_top_2')
// (2, 2, 'sp4_h_r_1')
// (2, 2, 'sp4_v_t_36')
// (2, 3, 'local_g2_2')
// (2, 3, 'lutff_1/in_1')
// (2, 3, 'lutff_2/out')
// (2, 3, 'sp4_v_b_36')
// (2, 4, 'neigh_op_bot_2')
// (2, 4, 'sp4_v_b_25')
// (2, 5, 'sp4_v_b_12')
// (2, 6, 'local_g0_1')
// (2, 6, 'lutff_2/in_1')
// (2, 6, 'sp4_v_b_1')
// (3, 2, 'neigh_op_tnl_2')
// (3, 2, 'sp4_h_r_12')
// (3, 3, 'neigh_op_lft_2')
// (3, 4, 'neigh_op_bnl_2')
// (4, 2, 'local_g2_1')
// (4, 2, 'lutff_5/in_0')
// (4, 2, 'sp4_h_r_25')
// (5, 2, 'sp4_h_r_36')
// (6, 2, 'sp4_h_l_36')

wire n53;
// (1, 2, 'neigh_op_tnr_3')
// (1, 3, 'local_g3_3')
// (1, 3, 'lutff_global/cen')
// (1, 3, 'neigh_op_rgt_3')
// (1, 4, 'neigh_op_bnr_3')
// (2, 2, 'neigh_op_top_3')
// (2, 3, 'local_g3_3')
// (2, 3, 'lutff_3/out')
// (2, 3, 'lutff_global/cen')
// (2, 4, 'neigh_op_bot_3')
// (3, 2, 'neigh_op_tnl_3')
// (3, 3, 'neigh_op_lft_3')
// (3, 4, 'neigh_op_bnl_3')

wire n54;
// (1, 2, 'neigh_op_tnr_4')
// (1, 3, 'neigh_op_rgt_4')
// (1, 4, 'neigh_op_bnr_4')
// (2, 2, 'neigh_op_top_4')
// (2, 3, 'local_g2_4')
// (2, 3, 'lutff_1/in_3')
// (2, 3, 'lutff_4/out')
// (2, 4, 'neigh_op_bot_4')
// (3, 2, 'neigh_op_tnl_4')
// (3, 3, 'neigh_op_lft_4')
// (3, 4, 'neigh_op_bnl_4')

wire n55;
// (1, 2, 'neigh_op_tnr_5')
// (1, 3, 'neigh_op_rgt_5')
// (1, 4, 'neigh_op_bnr_5')
// (2, 2, 'local_g0_5')
// (2, 2, 'lutff_1/in_2')
// (2, 2, 'neigh_op_top_5')
// (2, 3, 'lutff_5/out')
// (2, 3, 'sp4_r_v_b_43')
// (2, 4, 'neigh_op_bot_5')
// (2, 4, 'sp4_r_v_b_30')
// (2, 5, 'sp4_r_v_b_19')
// (2, 6, 'sp4_r_v_b_6')
// (3, 2, 'neigh_op_tnl_5')
// (3, 2, 'sp4_h_r_6')
// (3, 2, 'sp4_v_t_43')
// (3, 3, 'neigh_op_lft_5')
// (3, 3, 'sp4_v_b_43')
// (3, 4, 'neigh_op_bnl_5')
// (3, 4, 'sp4_v_b_30')
// (3, 5, 'sp4_v_b_19')
// (3, 6, 'sp4_v_b_6')
// (4, 2, 'local_g0_3')
// (4, 2, 'lutff_5/in_2')
// (4, 2, 'sp4_h_r_19')
// (5, 2, 'sp4_h_r_30')
// (6, 2, 'sp4_h_r_43')
// (7, 2, 'sp4_h_l_43')

reg n56 = 0;
// (1, 2, 'neigh_op_tnr_7')
// (1, 3, 'local_g2_7')
// (1, 3, 'lutff_0/in_1')
// (1, 3, 'lutff_4/in_3')
// (1, 3, 'neigh_op_rgt_7')
// (1, 4, 'neigh_op_bnr_7')
// (2, 2, 'neigh_op_top_7')
// (2, 3, 'local_g0_7')
// (2, 3, 'local_g1_7')
// (2, 3, 'lutff_0/in_3')
// (2, 3, 'lutff_2/in_3')
// (2, 3, 'lutff_5/in_3')
// (2, 3, 'lutff_6/in_3')
// (2, 3, 'lutff_7/in_3')
// (2, 3, 'lutff_7/out')
// (2, 4, 'neigh_op_bot_7')
// (3, 2, 'neigh_op_tnl_7')
// (3, 3, 'neigh_op_lft_7')
// (3, 4, 'neigh_op_bnl_7')

wire n57;
// (1, 3, 'lutff_1/cout')
// (1, 3, 'lutff_2/in_3')

wire n58;
// (1, 3, 'lutff_2/cout')
// (1, 3, 'lutff_3/in_3')

wire n59;
// (1, 3, 'neigh_op_tnr_7')
// (1, 4, 'neigh_op_rgt_7')
// (1, 5, 'neigh_op_bnr_7')
// (2, 0, 'span12_vert_21')
// (2, 1, 'sp12_v_b_21')
// (2, 2, 'sp12_v_b_18')
// (2, 2, 'sp4_r_v_b_39')
// (2, 3, 'local_g2_1')
// (2, 3, 'lutff_7/in_2')
// (2, 3, 'neigh_op_top_7')
// (2, 3, 'sp12_v_b_17')
// (2, 3, 'sp4_r_v_b_26')
// (2, 3, 'sp4_r_v_b_42')
// (2, 4, 'lutff_7/out')
// (2, 4, 'sp12_v_b_14')
// (2, 4, 'sp4_r_v_b_15')
// (2, 4, 'sp4_r_v_b_31')
// (2, 5, 'neigh_op_bot_7')
// (2, 5, 'sp12_v_b_13')
// (2, 5, 'sp4_r_v_b_18')
// (2, 5, 'sp4_r_v_b_2')
// (2, 6, 'sp12_v_b_10')
// (2, 6, 'sp4_r_v_b_7')
// (2, 7, 'sp12_v_b_9')
// (2, 8, 'sp12_v_b_6')
// (2, 9, 'sp12_v_b_5')
// (2, 10, 'sp12_v_b_2')
// (2, 11, 'sp12_v_b_1')
// (3, 1, 'sp4_v_t_39')
// (3, 2, 'sp4_v_b_39')
// (3, 2, 'sp4_v_t_42')
// (3, 3, 'neigh_op_tnl_7')
// (3, 3, 'sp4_v_b_26')
// (3, 3, 'sp4_v_b_42')
// (3, 4, 'neigh_op_lft_7')
// (3, 4, 'sp4_v_b_15')
// (3, 4, 'sp4_v_b_31')
// (3, 5, 'neigh_op_bnl_7')
// (3, 5, 'sp4_h_r_2')
// (3, 5, 'sp4_v_b_18')
// (3, 5, 'sp4_v_b_2')
// (3, 6, 'sp4_h_r_1')
// (3, 6, 'sp4_v_b_7')
// (4, 5, 'sp4_h_r_15')
// (4, 6, 'local_g1_4')
// (4, 6, 'lutff_2/in_3')
// (4, 6, 'sp4_h_r_12')
// (5, 5, 'sp4_h_r_26')
// (5, 6, 'local_g3_1')
// (5, 6, 'lutff_0/in_0')
// (5, 6, 'sp4_h_r_25')
// (6, 3, 'sp4_r_v_b_42')
// (6, 4, 'sp4_r_v_b_31')
// (6, 5, 'sp4_h_r_39')
// (6, 5, 'sp4_r_v_b_18')
// (6, 6, 'sp4_h_r_36')
// (6, 6, 'sp4_r_v_b_7')
// (7, 2, 'sp4_v_t_42')
// (7, 3, 'sp4_v_b_42')
// (7, 4, 'sp4_v_b_31')
// (7, 5, 'local_g0_2')
// (7, 5, 'lutff_3/in_3')
// (7, 5, 'sp4_h_l_39')
// (7, 5, 'sp4_h_r_10')
// (7, 5, 'sp4_v_b_18')
// (7, 6, 'local_g0_7')
// (7, 6, 'local_g1_7')
// (7, 6, 'lutff_0/in_0')
// (7, 6, 'lutff_5/in_0')
// (7, 6, 'sp4_h_l_36')
// (7, 6, 'sp4_v_b_7')
// (8, 5, 'local_g0_7')
// (8, 5, 'lutff_0/in_3')
// (8, 5, 'lutff_1/in_0')
// (8, 5, 'lutff_4/in_3')
// (8, 5, 'sp4_h_r_23')
// (9, 5, 'sp4_h_r_34')
// (10, 5, 'sp4_h_r_47')
// (11, 5, 'sp4_h_l_47')

reg n60 = 0;
// (1, 3, 'sp4_h_r_4')
// (2, 3, 'local_g0_1')
// (2, 3, 'lutff_4/in_1')
// (2, 3, 'lutff_7/in_0')
// (2, 3, 'sp4_h_r_17')
// (3, 2, 'neigh_op_tnr_5')
// (3, 3, 'neigh_op_rgt_5')
// (3, 3, 'sp4_h_r_28')
// (3, 4, 'neigh_op_bnr_5')
// (4, 1, 'sp4_r_v_b_35')
// (4, 2, 'neigh_op_top_5')
// (4, 2, 'sp4_r_v_b_22')
// (4, 3, 'local_g0_5')
// (4, 3, 'local_g1_5')
// (4, 3, 'lutff_0/in_3')
// (4, 3, 'lutff_2/in_3')
// (4, 3, 'lutff_5/in_1')
// (4, 3, 'lutff_5/out')
// (4, 3, 'sp4_h_r_41')
// (4, 3, 'sp4_r_v_b_11')
// (4, 4, 'neigh_op_bot_5')
// (5, 0, 'span4_vert_35')
// (5, 1, 'sp4_v_b_35')
// (5, 2, 'neigh_op_tnl_5')
// (5, 2, 'sp4_v_b_22')
// (5, 3, 'neigh_op_lft_5')
// (5, 3, 'sp4_h_l_41')
// (5, 3, 'sp4_v_b_11')
// (5, 4, 'neigh_op_bnl_5')

reg n61 = 0;
// (1, 4, 'neigh_op_tnr_2')
// (1, 5, 'neigh_op_rgt_2')
// (1, 6, 'neigh_op_bnr_2')
// (2, 4, 'neigh_op_top_2')
// (2, 5, 'local_g0_2')
// (2, 5, 'lutff_2/in_2')
// (2, 5, 'lutff_2/out')
// (2, 6, 'local_g0_2')
// (2, 6, 'local_g1_2')
// (2, 6, 'lutff_0/in_2')
// (2, 6, 'lutff_7/in_2')
// (2, 6, 'neigh_op_bot_2')
// (3, 4, 'neigh_op_tnl_2')
// (3, 5, 'neigh_op_lft_2')
// (3, 6, 'neigh_op_bnl_2')

reg n62 = 0;
// (1, 4, 'neigh_op_tnr_3')
// (1, 5, 'neigh_op_rgt_3')
// (1, 6, 'neigh_op_bnr_3')
// (2, 4, 'neigh_op_top_3')
// (2, 5, 'local_g0_3')
// (2, 5, 'lutff_3/in_2')
// (2, 5, 'lutff_3/out')
// (2, 6, 'local_g0_3')
// (2, 6, 'lutff_0/in_1')
// (2, 6, 'lutff_6/in_1')
// (2, 6, 'lutff_7/in_0')
// (2, 6, 'neigh_op_bot_3')
// (3, 4, 'neigh_op_tnl_3')
// (3, 5, 'neigh_op_lft_3')
// (3, 6, 'neigh_op_bnl_3')

reg n63 = 0;
// (1, 4, 'neigh_op_tnr_4')
// (1, 4, 'sp4_r_v_b_37')
// (1, 5, 'neigh_op_rgt_4')
// (1, 5, 'sp4_h_r_1')
// (1, 5, 'sp4_r_v_b_24')
// (1, 6, 'neigh_op_bnr_4')
// (1, 6, 'sp4_r_v_b_13')
// (1, 7, 'sp4_r_v_b_0')
// (2, 3, 'sp4_v_t_37')
// (2, 4, 'neigh_op_top_4')
// (2, 4, 'sp4_v_b_37')
// (2, 5, 'local_g0_4')
// (2, 5, 'lutff_4/in_2')
// (2, 5, 'lutff_4/out')
// (2, 5, 'sp12_h_r_0')
// (2, 5, 'sp4_h_r_12')
// (2, 5, 'sp4_v_b_24')
// (2, 6, 'local_g1_5')
// (2, 6, 'lutff_3/in_1')
// (2, 6, 'lutff_5/in_3')
// (2, 6, 'neigh_op_bot_4')
// (2, 6, 'sp4_v_b_13')
// (2, 7, 'sp4_v_b_0')
// (3, 4, 'neigh_op_tnl_4')
// (3, 5, 'neigh_op_lft_4')
// (3, 5, 'sp12_h_r_3')
// (3, 5, 'sp4_h_r_25')
// (3, 5, 'sp4_h_r_3')
// (3, 6, 'neigh_op_bnl_4')
// (4, 5, 'sp12_h_r_4')
// (4, 5, 'sp4_h_r_14')
// (4, 5, 'sp4_h_r_36')
// (4, 6, 'local_g2_4')
// (4, 6, 'lutff_0/in_2')
// (4, 6, 'lutff_4/in_0')
// (4, 6, 'sp4_r_v_b_36')
// (4, 7, 'sp4_r_v_b_25')
// (4, 8, 'sp4_r_v_b_12')
// (4, 9, 'sp4_r_v_b_1')
// (5, 5, 'sp12_h_r_7')
// (5, 5, 'sp4_h_l_36')
// (5, 5, 'sp4_h_r_27')
// (5, 5, 'sp4_h_r_5')
// (5, 5, 'sp4_v_t_36')
// (5, 6, 'sp4_v_b_36')
// (5, 7, 'sp4_v_b_25')
// (5, 8, 'sp4_v_b_12')
// (5, 9, 'sp4_v_b_1')
// (6, 5, 'sp12_h_r_8')
// (6, 5, 'sp4_h_r_16')
// (6, 5, 'sp4_h_r_38')
// (6, 6, 'sp4_r_v_b_38')
// (6, 7, 'sp4_r_v_b_27')
// (6, 8, 'sp4_r_v_b_14')
// (6, 9, 'sp4_r_v_b_3')
// (7, 5, 'local_g0_3')
// (7, 5, 'local_g3_5')
// (7, 5, 'lutff_0/in_0')
// (7, 5, 'lutff_4/in_1')
// (7, 5, 'lutff_7/in_1')
// (7, 5, 'sp12_h_r_11')
// (7, 5, 'sp4_h_l_38')
// (7, 5, 'sp4_h_r_29')
// (7, 5, 'sp4_v_t_38')
// (7, 6, 'local_g2_6')
// (7, 6, 'local_g3_6')
// (7, 6, 'lutff_3/in_3')
// (7, 6, 'lutff_4/in_3')
// (7, 6, 'sp4_v_b_38')
// (7, 7, 'sp4_v_b_27')
// (7, 8, 'sp4_v_b_14')
// (7, 9, 'sp4_v_b_3')
// (8, 5, 'sp12_h_r_12')
// (8, 5, 'sp4_h_r_40')
// (9, 5, 'sp12_h_r_15')
// (9, 5, 'sp4_h_l_40')
// (10, 5, 'sp12_h_r_16')
// (11, 5, 'sp12_h_r_19')
// (12, 5, 'sp12_h_r_20')
// (13, 5, 'span12_horz_20')

wire n64;
// (1, 5, 'neigh_op_tnr_0')
// (1, 6, 'neigh_op_rgt_0')
// (1, 7, 'neigh_op_bnr_0')
// (2, 5, 'neigh_op_top_0')
// (2, 6, 'local_g0_0')
// (2, 6, 'lutff_0/out')
// (2, 6, 'lutff_1/in_1')
// (2, 7, 'neigh_op_bot_0')
// (3, 5, 'neigh_op_tnl_0')
// (3, 6, 'neigh_op_lft_0')
// (3, 7, 'neigh_op_bnl_0')

wire n65;
// (1, 5, 'neigh_op_tnr_1')
// (1, 5, 'sp4_r_v_b_47')
// (1, 6, 'neigh_op_rgt_1')
// (1, 6, 'sp4_r_v_b_34')
// (1, 7, 'neigh_op_bnr_1')
// (1, 7, 'sp4_r_v_b_23')
// (1, 8, 'sp4_r_v_b_10')
// (2, 4, 'sp4_v_t_47')
// (2, 5, 'neigh_op_top_1')
// (2, 5, 'sp4_v_b_47')
// (2, 6, 'lutff_1/out')
// (2, 6, 'sp4_v_b_34')
// (2, 7, 'neigh_op_bot_1')
// (2, 7, 'sp4_v_b_23')
// (2, 8, 'local_g0_2')
// (2, 8, 'lutff_global/cen')
// (2, 8, 'sp4_v_b_10')
// (3, 5, 'neigh_op_tnl_1')
// (3, 6, 'neigh_op_lft_1')
// (3, 7, 'neigh_op_bnl_1')

wire n66;
// (1, 5, 'neigh_op_tnr_3')
// (1, 6, 'neigh_op_rgt_3')
// (1, 7, 'neigh_op_bnr_3')
// (2, 5, 'neigh_op_top_3')
// (2, 6, 'local_g1_3')
// (2, 6, 'lutff_2/in_2')
// (2, 6, 'lutff_3/out')
// (2, 7, 'neigh_op_bot_3')
// (3, 5, 'neigh_op_tnl_3')
// (3, 6, 'neigh_op_lft_3')
// (3, 7, 'neigh_op_bnl_3')

wire n67;
// (1, 5, 'neigh_op_tnr_5')
// (1, 6, 'neigh_op_rgt_5')
// (1, 7, 'neigh_op_bnr_5')
// (2, 5, 'neigh_op_top_5')
// (2, 6, 'local_g0_5')
// (2, 6, 'lutff_1/in_2')
// (2, 6, 'lutff_5/out')
// (2, 7, 'neigh_op_bot_5')
// (3, 5, 'neigh_op_tnl_5')
// (3, 6, 'neigh_op_lft_5')
// (3, 7, 'neigh_op_bnl_5')

reg n68 = 0;
// (1, 5, 'neigh_op_tnr_7')
// (1, 6, 'neigh_op_rgt_7')
// (1, 6, 'sp4_h_r_3')
// (1, 7, 'neigh_op_bnr_7')
// (2, 5, 'neigh_op_top_7')
// (2, 6, 'lutff_7/out')
// (2, 6, 'sp4_h_r_14')
// (2, 6, 'sp4_r_v_b_47')
// (2, 7, 'neigh_op_bot_7')
// (2, 7, 'sp4_r_v_b_34')
// (2, 8, 'sp4_r_v_b_23')
// (2, 9, 'sp4_r_v_b_10')
// (3, 5, 'neigh_op_tnl_7')
// (3, 5, 'sp4_v_t_47')
// (3, 6, 'neigh_op_lft_7')
// (3, 6, 'sp4_h_r_27')
// (3, 6, 'sp4_v_b_47')
// (3, 7, 'neigh_op_bnl_7')
// (3, 7, 'sp4_v_b_34')
// (3, 8, 'sp4_v_b_23')
// (3, 9, 'sp4_h_r_4')
// (3, 9, 'sp4_v_b_10')
// (3, 13, 'sp4_h_r_2')
// (4, 6, 'sp4_h_r_38')
// (4, 7, 'sp4_r_v_b_45')
// (4, 8, 'sp4_r_v_b_32')
// (4, 9, 'local_g0_1')
// (4, 9, 'lutff_3/in_2')
// (4, 9, 'sp4_h_r_17')
// (4, 9, 'sp4_r_v_b_21')
// (4, 10, 'sp4_r_v_b_8')
// (4, 11, 'sp4_r_v_b_46')
// (4, 12, 'sp4_r_v_b_35')
// (4, 13, 'sp4_h_r_15')
// (4, 13, 'sp4_r_v_b_22')
// (4, 14, 'sp4_r_v_b_11')
// (5, 6, 'sp4_h_l_38')
// (5, 6, 'sp4_v_t_45')
// (5, 7, 'sp4_v_b_45')
// (5, 8, 'sp4_v_b_32')
// (5, 9, 'local_g2_4')
// (5, 9, 'lutff_7/in_3')
// (5, 9, 'sp4_h_r_28')
// (5, 9, 'sp4_v_b_21')
// (5, 10, 'local_g0_0')
// (5, 10, 'lutff_1/in_1')
// (5, 10, 'sp4_h_r_7')
// (5, 10, 'sp4_h_r_8')
// (5, 10, 'sp4_v_b_8')
// (5, 10, 'sp4_v_t_46')
// (5, 11, 'local_g2_6')
// (5, 11, 'local_g3_6')
// (5, 11, 'lutff_0/in_2')
// (5, 11, 'lutff_5/in_3')
// (5, 11, 'lutff_7/in_2')
// (5, 11, 'sp4_v_b_46')
// (5, 12, 'sp4_v_b_35')
// (5, 13, 'local_g2_2')
// (5, 13, 'local_g3_2')
// (5, 13, 'lutff_0/in_2')
// (5, 13, 'lutff_1/in_2')
// (5, 13, 'lutff_2/in_1')
// (5, 13, 'sp4_h_r_26')
// (5, 13, 'sp4_v_b_22')
// (5, 14, 'local_g0_3')
// (5, 14, 'local_g1_3')
// (5, 14, 'lutff_4/in_2')
// (5, 14, 'lutff_6/in_3')
// (5, 14, 'sp4_v_b_11')
// (6, 9, 'local_g2_1')
// (6, 9, 'local_g3_1')
// (6, 9, 'lutff_2/in_2')
// (6, 9, 'lutff_4/in_1')
// (6, 9, 'sp4_h_r_41')
// (6, 10, 'sp4_h_r_18')
// (6, 10, 'sp4_h_r_21')
// (6, 10, 'sp4_r_v_b_41')
// (6, 10, 'sp4_r_v_b_44')
// (6, 11, 'local_g0_2')
// (6, 11, 'lutff_2/in_2')
// (6, 11, 'sp4_r_v_b_28')
// (6, 11, 'sp4_r_v_b_33')
// (6, 12, 'local_g3_1')
// (6, 12, 'local_g3_4')
// (6, 12, 'lutff_0/in_1')
// (6, 12, 'lutff_2/in_2')
// (6, 12, 'lutff_3/in_1')
// (6, 12, 'lutff_6/in_3')
// (6, 12, 'sp4_r_v_b_17')
// (6, 12, 'sp4_r_v_b_20')
// (6, 13, 'local_g2_1')
// (6, 13, 'lutff_6/in_3')
// (6, 13, 'lutff_7/in_2')
// (6, 13, 'sp4_h_r_39')
// (6, 13, 'sp4_r_v_b_4')
// (6, 13, 'sp4_r_v_b_9')
// (6, 14, 'sp4_r_v_b_40')
// (6, 15, 'sp4_r_v_b_29')
// (6, 16, 'sp4_r_v_b_16')
// (7, 9, 'sp4_h_l_41')
// (7, 9, 'sp4_v_t_41')
// (7, 9, 'sp4_v_t_44')
// (7, 10, 'local_g2_4')
// (7, 10, 'local_g3_4')
// (7, 10, 'lutff_2/in_1')
// (7, 10, 'lutff_3/in_2')
// (7, 10, 'lutff_7/in_3')
// (7, 10, 'sp4_h_r_31')
// (7, 10, 'sp4_h_r_32')
// (7, 10, 'sp4_v_b_41')
// (7, 10, 'sp4_v_b_44')
// (7, 11, 'local_g2_1')
// (7, 11, 'lutff_2/in_1')
// (7, 11, 'sp4_v_b_28')
// (7, 11, 'sp4_v_b_33')
// (7, 12, 'local_g0_4')
// (7, 12, 'lutff_2/in_2')
// (7, 12, 'sp4_v_b_17')
// (7, 12, 'sp4_v_b_20')
// (7, 13, 'local_g0_1')
// (7, 13, 'lutff_3/in_2')
// (7, 13, 'sp4_h_l_39')
// (7, 13, 'sp4_v_b_4')
// (7, 13, 'sp4_v_b_9')
// (7, 13, 'sp4_v_t_40')
// (7, 14, 'local_g2_0')
// (7, 14, 'lutff_0/in_2')
// (7, 14, 'lutff_1/in_1')
// (7, 14, 'lutff_2/in_2')
// (7, 14, 'lutff_5/in_3')
// (7, 14, 'sp4_v_b_40')
// (7, 15, 'sp4_v_b_29')
// (7, 16, 'sp4_v_b_16')
// (7, 17, 'span4_vert_5')
// (8, 10, 'sp4_h_r_42')
// (8, 10, 'sp4_h_r_45')
// (8, 11, 'local_g2_4')
// (8, 11, 'local_g2_5')
// (8, 11, 'lutff_0/in_2')
// (8, 11, 'lutff_7/in_2')
// (8, 11, 'sp4_r_v_b_36')
// (8, 11, 'sp4_r_v_b_37')
// (8, 11, 'sp4_r_v_b_45')
// (8, 12, 'local_g0_3')
// (8, 12, 'lutff_2/in_3')
// (8, 12, 'sp4_r_v_b_24')
// (8, 12, 'sp4_r_v_b_25')
// (8, 12, 'sp4_r_v_b_32')
// (8, 13, 'sp4_r_v_b_12')
// (8, 13, 'sp4_r_v_b_13')
// (8, 13, 'sp4_r_v_b_21')
// (8, 14, 'sp4_r_v_b_0')
// (8, 14, 'sp4_r_v_b_1')
// (8, 14, 'sp4_r_v_b_8')
// (9, 10, 'sp4_h_l_42')
// (9, 10, 'sp4_h_l_45')
// (9, 10, 'sp4_v_t_36')
// (9, 10, 'sp4_v_t_37')
// (9, 10, 'sp4_v_t_45')
// (9, 11, 'sp4_v_b_36')
// (9, 11, 'sp4_v_b_37')
// (9, 11, 'sp4_v_b_45')
// (9, 12, 'sp4_v_b_24')
// (9, 12, 'sp4_v_b_25')
// (9, 12, 'sp4_v_b_32')
// (9, 13, 'sp4_v_b_12')
// (9, 13, 'sp4_v_b_13')
// (9, 13, 'sp4_v_b_21')
// (9, 14, 'sp4_v_b_0')
// (9, 14, 'sp4_v_b_1')
// (9, 14, 'sp4_v_b_8')

wire n69;
// (1, 5, 'sp12_h_r_0')
// (2, 5, 'sp12_h_r_3')
// (3, 5, 'sp12_h_r_4')
// (4, 4, 'neigh_op_tnr_0')
// (4, 5, 'neigh_op_rgt_0')
// (4, 5, 'sp12_h_r_7')
// (4, 6, 'neigh_op_bnr_0')
// (5, 4, 'neigh_op_top_0')
// (5, 5, 'lutff_0/out')
// (5, 5, 'sp12_h_r_8')
// (5, 6, 'neigh_op_bot_0')
// (6, 4, 'neigh_op_tnl_0')
// (6, 5, 'local_g1_0')
// (6, 5, 'local_g1_3')
// (6, 5, 'lutff_5/in_0')
// (6, 5, 'lutff_6/in_2')
// (6, 5, 'neigh_op_lft_0')
// (6, 5, 'sp12_h_r_11')
// (6, 6, 'neigh_op_bnl_0')
// (7, 5, 'sp12_h_r_12')
// (8, 5, 'sp12_h_r_15')
// (9, 5, 'sp12_h_r_16')
// (10, 5, 'sp12_h_r_19')
// (11, 5, 'sp12_h_r_20')
// (12, 5, 'sp12_h_r_23')
// (13, 5, 'span12_horz_23')

reg n70 = 0;
// (1, 6, 'neigh_op_tnr_7')
// (1, 7, 'neigh_op_rgt_7')
// (1, 7, 'sp4_r_v_b_46')
// (1, 8, 'neigh_op_bnr_7')
// (1, 8, 'sp4_r_v_b_35')
// (1, 9, 'sp4_r_v_b_22')
// (1, 10, 'sp4_r_v_b_11')
// (2, 6, 'neigh_op_top_7')
// (2, 6, 'sp4_r_v_b_42')
// (2, 6, 'sp4_v_t_46')
// (2, 7, 'lutff_7/out')
// (2, 7, 'sp4_r_v_b_31')
// (2, 7, 'sp4_v_b_46')
// (2, 8, 'neigh_op_bot_7')
// (2, 8, 'sp4_r_v_b_18')
// (2, 8, 'sp4_v_b_35')
// (2, 9, 'sp4_r_v_b_7')
// (2, 9, 'sp4_v_b_22')
// (2, 10, 'sp4_h_r_11')
// (2, 10, 'sp4_v_b_11')
// (3, 5, 'sp4_h_r_7')
// (3, 5, 'sp4_v_t_42')
// (3, 6, 'neigh_op_tnl_7')
// (3, 6, 'sp4_v_b_42')
// (3, 7, 'neigh_op_lft_7')
// (3, 7, 'sp4_v_b_31')
// (3, 8, 'neigh_op_bnl_7')
// (3, 8, 'sp4_v_b_18')
// (3, 9, 'sp4_v_b_7')
// (3, 10, 'sp4_h_r_22')
// (3, 13, 'sp4_h_r_0')
// (4, 5, 'sp4_h_r_18')
// (4, 10, 'sp4_h_r_35')
// (4, 13, 'sp4_h_r_13')
// (5, 5, 'sp4_h_r_31')
// (5, 10, 'sp4_h_r_46')
// (5, 11, 'sp4_r_v_b_46')
// (5, 12, 'sp4_r_v_b_35')
// (5, 13, 'sp4_h_r_24')
// (5, 13, 'sp4_r_v_b_22')
// (5, 14, 'sp4_r_v_b_11')
// (6, 5, 'sp4_h_r_42')
// (6, 6, 'sp4_r_v_b_42')
// (6, 7, 'sp4_r_v_b_31')
// (6, 8, 'sp4_r_v_b_18')
// (6, 9, 'sp4_r_v_b_7')
// (6, 10, 'sp4_h_l_46')
// (6, 10, 'sp4_h_r_11')
// (6, 10, 'sp4_r_v_b_42')
// (6, 10, 'sp4_v_t_46')
// (6, 11, 'sp4_r_v_b_31')
// (6, 11, 'sp4_v_b_46')
// (6, 12, 'sp4_r_v_b_18')
// (6, 12, 'sp4_v_b_35')
// (6, 13, 'sp4_h_r_37')
// (6, 13, 'sp4_r_v_b_7')
// (6, 13, 'sp4_v_b_22')
// (6, 14, 'local_g0_3')
// (6, 14, 'lutff_6/in_3')
// (6, 14, 'sp4_v_b_11')
// (7, 5, 'sp4_h_l_42')
// (7, 5, 'sp4_h_r_0')
// (7, 5, 'sp4_v_t_42')
// (7, 6, 'sp4_v_b_42')
// (7, 7, 'sp4_v_b_31')
// (7, 8, 'sp4_v_b_18')
// (7, 9, 'local_g0_7')
// (7, 9, 'lutff_0/in_3')
// (7, 9, 'sp4_h_r_0')
// (7, 9, 'sp4_v_b_7')
// (7, 9, 'sp4_v_t_42')
// (7, 10, 'local_g0_6')
// (7, 10, 'lutff_1/in_3')
// (7, 10, 'sp4_h_r_22')
// (7, 10, 'sp4_v_b_42')
// (7, 11, 'local_g2_7')
// (7, 11, 'lutff_0/in_3')
// (7, 11, 'sp4_v_b_31')
// (7, 12, 'sp4_v_b_18')
// (7, 13, 'sp4_h_l_37')
// (7, 13, 'sp4_h_r_0')
// (7, 13, 'sp4_h_r_7')
// (7, 13, 'sp4_v_b_7')
// (8, 5, 'sp4_h_r_13')
// (8, 6, 'sp4_r_v_b_40')
// (8, 7, 'sp4_r_v_b_29')
// (8, 8, 'sp4_r_v_b_16')
// (8, 9, 'local_g1_5')
// (8, 9, 'lutff_5/in_3')
// (8, 9, 'lutff_7/in_3')
// (8, 9, 'sp4_h_r_13')
// (8, 9, 'sp4_r_v_b_5')
// (8, 10, 'local_g2_3')
// (8, 10, 'local_g3_3')
// (8, 10, 'lutff_3/in_3')
// (8, 10, 'lutff_4/in_3')
// (8, 10, 'sp4_h_r_35')
// (8, 10, 'sp4_r_v_b_36')
// (8, 10, 'sp4_r_v_b_37')
// (8, 11, 'local_g1_0')
// (8, 11, 'lutff_4/in_3')
// (8, 11, 'lutff_6/in_3')
// (8, 11, 'sp4_r_v_b_24')
// (8, 11, 'sp4_r_v_b_25')
// (8, 12, 'local_g2_4')
// (8, 12, 'lutff_1/in_3')
// (8, 12, 'sp4_r_v_b_12')
// (8, 12, 'sp4_r_v_b_13')
// (8, 13, 'local_g0_2')
// (8, 13, 'local_g0_5')
// (8, 13, 'lutff_0/in_3')
// (8, 13, 'lutff_2/in_3')
// (8, 13, 'lutff_7/in_3')
// (8, 13, 'sp4_h_r_13')
// (8, 13, 'sp4_h_r_18')
// (8, 13, 'sp4_r_v_b_0')
// (8, 13, 'sp4_r_v_b_1')
// (9, 5, 'sp4_h_r_24')
// (9, 5, 'sp4_v_t_40')
// (9, 6, 'sp4_v_b_40')
// (9, 7, 'sp4_r_v_b_38')
// (9, 7, 'sp4_r_v_b_46')
// (9, 7, 'sp4_v_b_29')
// (9, 8, 'sp4_r_v_b_27')
// (9, 8, 'sp4_r_v_b_35')
// (9, 8, 'sp4_v_b_16')
// (9, 9, 'local_g2_6')
// (9, 9, 'local_g3_6')
// (9, 9, 'lutff_0/in_3')
// (9, 9, 'lutff_1/in_3')
// (9, 9, 'lutff_3/in_3')
// (9, 9, 'lutff_6/in_3')
// (9, 9, 'sp4_h_r_0')
// (9, 9, 'sp4_h_r_24')
// (9, 9, 'sp4_r_v_b_14')
// (9, 9, 'sp4_r_v_b_22')
// (9, 9, 'sp4_v_b_5')
// (9, 9, 'sp4_v_t_36')
// (9, 9, 'sp4_v_t_37')
// (9, 10, 'sp4_h_r_46')
// (9, 10, 'sp4_r_v_b_11')
// (9, 10, 'sp4_r_v_b_3')
// (9, 10, 'sp4_v_b_36')
// (9, 10, 'sp4_v_b_37')
// (9, 11, 'sp4_r_v_b_41')
// (9, 11, 'sp4_r_v_b_42')
// (9, 11, 'sp4_v_b_24')
// (9, 11, 'sp4_v_b_25')
// (9, 12, 'local_g0_4')
// (9, 12, 'local_g0_7')
// (9, 12, 'lutff_0/in_3')
// (9, 12, 'lutff_2/in_3')
// (9, 12, 'lutff_3/in_3')
// (9, 12, 'lutff_4/in_3')
// (9, 12, 'lutff_5/in_3')
// (9, 12, 'sp4_r_v_b_28')
// (9, 12, 'sp4_r_v_b_31')
// (9, 12, 'sp4_v_b_12')
// (9, 12, 'sp4_v_b_13')
// (9, 13, 'sp4_h_r_24')
// (9, 13, 'sp4_h_r_31')
// (9, 13, 'sp4_r_v_b_17')
// (9, 13, 'sp4_r_v_b_18')
// (9, 13, 'sp4_v_b_0')
// (9, 13, 'sp4_v_b_1')
// (9, 14, 'sp4_r_v_b_4')
// (9, 14, 'sp4_r_v_b_7')
// (10, 5, 'sp4_h_r_37')
// (10, 6, 'sp4_r_v_b_40')
// (10, 6, 'sp4_v_t_38')
// (10, 6, 'sp4_v_t_46')
// (10, 7, 'sp4_r_v_b_29')
// (10, 7, 'sp4_v_b_38')
// (10, 7, 'sp4_v_b_46')
// (10, 8, 'sp4_r_v_b_16')
// (10, 8, 'sp4_v_b_27')
// (10, 8, 'sp4_v_b_35')
// (10, 9, 'sp4_h_r_13')
// (10, 9, 'sp4_h_r_37')
// (10, 9, 'sp4_r_v_b_5')
// (10, 9, 'sp4_v_b_14')
// (10, 9, 'sp4_v_b_22')
// (10, 10, 'sp4_h_l_46')
// (10, 10, 'sp4_v_b_11')
// (10, 10, 'sp4_v_b_3')
// (10, 10, 'sp4_v_t_41')
// (10, 10, 'sp4_v_t_42')
// (10, 11, 'sp4_v_b_41')
// (10, 11, 'sp4_v_b_42')
// (10, 12, 'sp4_v_b_28')
// (10, 12, 'sp4_v_b_31')
// (10, 13, 'sp4_h_r_37')
// (10, 13, 'sp4_h_r_42')
// (10, 13, 'sp4_v_b_17')
// (10, 13, 'sp4_v_b_18')
// (10, 14, 'sp4_v_b_4')
// (10, 14, 'sp4_v_b_7')
// (11, 5, 'sp4_h_l_37')
// (11, 5, 'sp4_v_t_40')
// (11, 6, 'sp4_v_b_40')
// (11, 7, 'sp4_v_b_29')
// (11, 8, 'sp4_v_b_16')
// (11, 9, 'local_g1_5')
// (11, 9, 'lutff_3/in_3')
// (11, 9, 'lutff_7/in_3')
// (11, 9, 'sp4_h_l_37')
// (11, 9, 'sp4_h_r_0')
// (11, 9, 'sp4_h_r_24')
// (11, 9, 'sp4_v_b_5')
// (11, 13, 'sp4_h_l_37')
// (11, 13, 'sp4_h_l_42')
// (12, 9, 'sp4_h_r_13')
// (12, 9, 'sp4_h_r_37')
// (13, 9, 'span4_horz_13')
// (13, 9, 'span4_horz_37')

wire n71;
// (1, 6, 'sp4_h_r_10')
// (2, 6, 'sp4_h_r_23')
// (3, 6, 'sp4_h_r_34')
// (4, 6, 'sp4_h_r_47')
// (4, 7, 'sp4_r_v_b_47')
// (4, 8, 'sp4_r_v_b_34')
// (4, 9, 'sp4_r_v_b_23')
// (4, 10, 'sp4_r_v_b_10')
// (5, 6, 'sp4_h_l_47')
// (5, 6, 'sp4_h_r_2')
// (5, 6, 'sp4_v_t_47')
// (5, 7, 'local_g2_7')
// (5, 7, 'lutff_5/in_0')
// (5, 7, 'sp4_v_b_47')
// (5, 8, 'sp4_v_b_34')
// (5, 9, 'sp4_v_b_23')
// (5, 10, 'sp4_v_b_10')
// (6, 5, 'neigh_op_tnr_5')
// (6, 6, 'neigh_op_rgt_5')
// (6, 6, 'sp4_h_r_15')
// (6, 7, 'neigh_op_bnr_5')
// (7, 5, 'neigh_op_top_5')
// (7, 6, 'lutff_5/out')
// (7, 6, 'sp4_h_r_10')
// (7, 6, 'sp4_h_r_26')
// (7, 7, 'neigh_op_bot_5')
// (8, 5, 'neigh_op_tnl_5')
// (8, 6, 'neigh_op_lft_5')
// (8, 6, 'sp4_h_r_23')
// (8, 6, 'sp4_h_r_39')
// (8, 7, 'neigh_op_bnl_5')
// (9, 6, 'sp4_h_l_39')
// (9, 6, 'sp4_h_r_34')
// (10, 6, 'sp4_h_r_47')
// (10, 7, 'sp4_r_v_b_47')
// (10, 8, 'sp4_r_v_b_34')
// (10, 9, 'sp4_r_v_b_23')
// (10, 10, 'sp4_r_v_b_10')
// (11, 6, 'sp4_h_l_47')
// (11, 6, 'sp4_v_t_47')
// (11, 7, 'local_g2_7')
// (11, 7, 'lutff_1/in_2')
// (11, 7, 'lutff_7/in_2')
// (11, 7, 'sp4_v_b_47')
// (11, 8, 'sp4_v_b_34')
// (11, 9, 'sp4_v_b_23')
// (11, 10, 'sp4_v_b_10')

wire n72;
// (1, 6, 'sp4_h_r_11')
// (1, 6, 'sp4_v_t_40')
// (1, 7, 'local_g2_0')
// (1, 7, 'lutff_4/in_0')
// (1, 7, 'sp4_v_b_40')
// (1, 8, 'sp4_v_b_29')
// (1, 9, 'sp4_v_b_16')
// (1, 10, 'sp4_v_b_5')
// (2, 6, 'sp4_h_r_22')
// (3, 6, 'sp4_h_r_35')
// (4, 6, 'sp4_h_r_46')
// (4, 7, 'sp4_r_v_b_39')
// (4, 8, 'sp4_r_v_b_26')
// (4, 9, 'sp4_r_v_b_15')
// (4, 10, 'local_g1_2')
// (4, 10, 'lutff_7/in_2')
// (4, 10, 'sp4_r_v_b_2')
// (5, 6, 'sp4_h_l_46')
// (5, 6, 'sp4_h_r_8')
// (5, 6, 'sp4_v_t_39')
// (5, 7, 'sp4_v_b_39')
// (5, 8, 'sp4_v_b_26')
// (5, 9, 'sp4_v_b_15')
// (5, 10, 'sp4_h_r_2')
// (5, 10, 'sp4_v_b_2')
// (6, 5, 'neigh_op_tnr_0')
// (6, 6, 'neigh_op_rgt_0')
// (6, 6, 'sp4_h_r_21')
// (6, 7, 'neigh_op_bnr_0')
// (6, 10, 'sp4_h_r_15')
// (7, 5, 'neigh_op_top_0')
// (7, 6, 'lutff_0/out')
// (7, 6, 'sp4_h_r_32')
// (7, 7, 'neigh_op_bot_0')
// (7, 10, 'sp4_h_r_26')
// (8, 5, 'neigh_op_tnl_0')
// (8, 6, 'neigh_op_lft_0')
// (8, 6, 'sp4_h_r_45')
// (8, 7, 'neigh_op_bnl_0')
// (8, 10, 'local_g2_7')
// (8, 10, 'lutff_5/in_2')
// (8, 10, 'sp4_h_r_39')
// (9, 6, 'sp4_h_l_45')
// (9, 10, 'sp4_h_l_39')

wire n73;
// (1, 7, 'sp4_h_r_10')
// (2, 7, 'local_g0_7')
// (2, 7, 'lutff_7/in_0')
// (2, 7, 'sp4_h_r_23')
// (3, 5, 'neigh_op_tnr_3')
// (3, 6, 'neigh_op_rgt_3')
// (3, 7, 'neigh_op_bnr_3')
// (3, 7, 'sp4_h_r_34')
// (4, 4, 'sp4_r_v_b_47')
// (4, 5, 'neigh_op_top_3')
// (4, 5, 'sp12_v_t_22')
// (4, 5, 'sp4_r_v_b_34')
// (4, 6, 'lutff_3/out')
// (4, 6, 'sp12_v_b_22')
// (4, 6, 'sp4_r_v_b_23')
// (4, 7, 'neigh_op_bot_3')
// (4, 7, 'sp12_v_b_21')
// (4, 7, 'sp4_h_r_47')
// (4, 7, 'sp4_r_v_b_10')
// (4, 8, 'local_g2_2')
// (4, 8, 'lutff_3/in_3')
// (4, 8, 'sp12_v_b_18')
// (4, 9, 'sp12_v_b_17')
// (4, 10, 'sp12_v_b_14')
// (4, 11, 'sp12_v_b_13')
// (4, 12, 'sp12_v_b_10')
// (4, 13, 'sp12_v_b_9')
// (4, 14, 'sp12_v_b_6')
// (4, 15, 'sp12_v_b_5')
// (4, 16, 'sp12_v_b_2')
// (4, 17, 'span12_vert_1')
// (5, 3, 'sp4_v_t_47')
// (5, 4, 'sp4_v_b_47')
// (5, 5, 'neigh_op_tnl_3')
// (5, 5, 'sp4_v_b_34')
// (5, 6, 'neigh_op_lft_3')
// (5, 6, 'sp4_v_b_23')
// (5, 7, 'neigh_op_bnl_3')
// (5, 7, 'sp4_h_l_47')
// (5, 7, 'sp4_v_b_10')

reg n74 = 0;
// (1, 7, 'sp4_r_v_b_38')
// (1, 8, 'neigh_op_tnr_7')
// (1, 8, 'sp4_r_v_b_27')
// (1, 9, 'neigh_op_rgt_7')
// (1, 9, 'sp4_r_v_b_14')
// (1, 10, 'neigh_op_bnr_7')
// (1, 10, 'sp4_r_v_b_3')
// (2, 6, 'sp4_v_t_38')
// (2, 7, 'sp4_v_b_38')
// (2, 8, 'neigh_op_top_7')
// (2, 8, 'sp4_v_b_27')
// (2, 9, 'lutff_7/out')
// (2, 9, 'sp4_v_b_14')
// (2, 10, 'local_g1_3')
// (2, 10, 'lutff_6/in_0')
// (2, 10, 'neigh_op_bot_7')
// (2, 10, 'sp4_v_b_3')
// (3, 8, 'neigh_op_tnl_7')
// (3, 9, 'neigh_op_lft_7')
// (3, 10, 'neigh_op_bnl_7')

reg n75 = 0;
// (1, 8, 'neigh_op_tnr_0')
// (1, 9, 'neigh_op_rgt_0')
// (1, 9, 'sp4_h_r_5')
// (1, 10, 'neigh_op_bnr_0')
// (2, 8, 'neigh_op_top_0')
// (2, 9, 'lutff_0/out')
// (2, 9, 'sp4_h_r_16')
// (2, 10, 'neigh_op_bot_0')
// (3, 8, 'neigh_op_tnl_0')
// (3, 9, 'neigh_op_lft_0')
// (3, 9, 'sp4_h_r_29')
// (3, 10, 'neigh_op_bnl_0')
// (4, 9, 'local_g2_0')
// (4, 9, 'lutff_4/in_0')
// (4, 9, 'sp4_h_r_40')
// (5, 9, 'sp4_h_l_40')

reg n76 = 0;
// (1, 8, 'neigh_op_tnr_2')
// (1, 9, 'neigh_op_rgt_2')
// (1, 10, 'neigh_op_bnr_2')
// (2, 8, 'neigh_op_top_2')
// (2, 9, 'local_g1_2')
// (2, 9, 'lutff_2/out')
// (2, 9, 'lutff_7/in_0')
// (2, 10, 'neigh_op_bot_2')
// (3, 8, 'neigh_op_tnl_2')
// (3, 9, 'neigh_op_lft_2')
// (3, 10, 'neigh_op_bnl_2')

reg n77 = 0;
// (1, 8, 'sp4_r_v_b_40')
// (1, 9, 'sp4_r_v_b_29')
// (1, 10, 'sp4_r_v_b_16')
// (1, 11, 'sp4_r_v_b_5')
// (2, 7, 'sp4_v_t_40')
// (2, 8, 'sp4_v_b_40')
// (2, 9, 'sp4_v_b_29')
// (2, 10, 'local_g0_0')
// (2, 10, 'lutff_4/in_0')
// (2, 10, 'sp4_v_b_16')
// (2, 11, 'sp4_h_r_0')
// (2, 11, 'sp4_v_b_5')
// (3, 10, 'neigh_op_tnr_4')
// (3, 11, 'neigh_op_rgt_4')
// (3, 11, 'sp4_h_r_13')
// (3, 12, 'neigh_op_bnr_4')
// (4, 10, 'neigh_op_top_4')
// (4, 11, 'lutff_4/out')
// (4, 11, 'sp4_h_r_24')
// (4, 12, 'neigh_op_bot_4')
// (5, 10, 'neigh_op_tnl_4')
// (5, 11, 'neigh_op_lft_4')
// (5, 11, 'sp4_h_r_37')
// (5, 12, 'neigh_op_bnl_4')
// (6, 11, 'sp4_h_l_37')

reg n78 = 0;
// (1, 9, 'neigh_op_tnr_1')
// (1, 10, 'neigh_op_rgt_1')
// (1, 11, 'neigh_op_bnr_1')
// (2, 9, 'neigh_op_top_1')
// (2, 9, 'sp4_r_v_b_46')
// (2, 10, 'lutff_1/out')
// (2, 10, 'sp4_r_v_b_35')
// (2, 11, 'neigh_op_bot_1')
// (2, 11, 'sp4_r_v_b_22')
// (2, 12, 'sp4_r_v_b_11')
// (3, 8, 'sp4_h_r_11')
// (3, 8, 'sp4_v_t_46')
// (3, 9, 'neigh_op_tnl_1')
// (3, 9, 'sp4_v_b_46')
// (3, 10, 'neigh_op_lft_1')
// (3, 10, 'sp4_v_b_35')
// (3, 11, 'neigh_op_bnl_1')
// (3, 11, 'sp4_v_b_22')
// (3, 12, 'sp4_v_b_11')
// (4, 8, 'local_g0_6')
// (4, 8, 'lutff_2/in_0')
// (4, 8, 'sp4_h_r_22')
// (5, 8, 'sp4_h_r_35')
// (6, 8, 'sp4_h_r_46')
// (7, 8, 'sp4_h_l_46')

reg n79 = 0;
// (1, 9, 'neigh_op_tnr_2')
// (1, 10, 'neigh_op_rgt_2')
// (1, 11, 'neigh_op_bnr_2')
// (2, 9, 'neigh_op_top_2')
// (2, 10, 'local_g0_2')
// (2, 10, 'lutff_0/in_0')
// (2, 10, 'lutff_2/out')
// (2, 11, 'neigh_op_bot_2')
// (3, 9, 'neigh_op_tnl_2')
// (3, 10, 'neigh_op_lft_2')
// (3, 11, 'neigh_op_bnl_2')

reg n80 = 0;
// (1, 9, 'neigh_op_tnr_4')
// (1, 10, 'neigh_op_rgt_4')
// (1, 11, 'neigh_op_bnr_4')
// (2, 9, 'neigh_op_top_4')
// (2, 10, 'local_g1_4')
// (2, 10, 'lutff_1/in_0')
// (2, 10, 'lutff_4/out')
// (2, 11, 'neigh_op_bot_4')
// (3, 9, 'neigh_op_tnl_4')
// (3, 10, 'neigh_op_lft_4')
// (3, 11, 'neigh_op_bnl_4')

reg n81 = 0;
// (1, 9, 'neigh_op_tnr_6')
// (1, 10, 'neigh_op_rgt_6')
// (1, 11, 'neigh_op_bnr_6')
// (2, 9, 'neigh_op_top_6')
// (2, 10, 'local_g1_6')
// (2, 10, 'lutff_6/out')
// (2, 10, 'lutff_7/in_0')
// (2, 11, 'neigh_op_bot_6')
// (3, 9, 'neigh_op_tnl_6')
// (3, 10, 'neigh_op_lft_6')
// (3, 11, 'neigh_op_bnl_6')

reg n82 = 0;
// (1, 9, 'neigh_op_tnr_7')
// (1, 10, 'neigh_op_rgt_7')
// (1, 11, 'neigh_op_bnr_7')
// (2, 9, 'neigh_op_top_7')
// (2, 10, 'local_g1_7')
// (2, 10, 'lutff_2/in_0')
// (2, 10, 'lutff_7/out')
// (2, 11, 'neigh_op_bot_7')
// (3, 9, 'neigh_op_tnl_7')
// (3, 10, 'neigh_op_lft_7')
// (3, 11, 'neigh_op_bnl_7')

reg n83 = 0;
// (1, 9, 'sp12_h_r_0')
// (2, 9, 'sp12_h_r_3')
// (3, 9, 'sp12_h_r_4')
// (4, 9, 'sp12_h_r_7')
// (5, 9, 'sp12_h_r_8')
// (6, 9, 'sp12_h_r_11')
// (7, 9, 'sp12_h_r_12')
// (8, 9, 'sp12_h_r_15')
// (9, 9, 'local_g0_0')
// (9, 9, 'lutff_0/in_2')
// (9, 9, 'sp12_h_r_16')
// (10, 8, 'neigh_op_tnr_6')
// (10, 9, 'neigh_op_rgt_6')
// (10, 9, 'sp12_h_r_19')
// (10, 10, 'neigh_op_bnr_6')
// (11, 8, 'neigh_op_top_6')
// (11, 9, 'local_g0_6')
// (11, 9, 'lutff_1/in_1')
// (11, 9, 'lutff_6/out')
// (11, 9, 'sp12_h_r_20')
// (11, 10, 'neigh_op_bot_6')
// (12, 8, 'neigh_op_tnl_6')
// (12, 9, 'neigh_op_lft_6')
// (12, 9, 'sp12_h_r_23')
// (12, 10, 'neigh_op_bnl_6')
// (13, 9, 'span12_horz_23')

reg n84 = 0;
// (1, 9, 'sp4_h_r_11')
// (2, 9, 'local_g1_6')
// (2, 9, 'lutff_3/in_0')
// (2, 9, 'sp4_h_r_22')
// (3, 8, 'neigh_op_tnr_7')
// (3, 9, 'neigh_op_rgt_7')
// (3, 9, 'sp4_h_r_35')
// (3, 10, 'neigh_op_bnr_7')
// (4, 8, 'neigh_op_top_7')
// (4, 9, 'lutff_7/out')
// (4, 9, 'sp4_h_r_46')
// (4, 10, 'neigh_op_bot_7')
// (5, 8, 'neigh_op_tnl_7')
// (5, 9, 'neigh_op_lft_7')
// (5, 9, 'sp4_h_l_46')
// (5, 10, 'neigh_op_bnl_7')

reg n85 = 0;
// (1, 10, 'neigh_op_tnr_4')
// (1, 11, 'neigh_op_rgt_4')
// (1, 12, 'neigh_op_bnr_4')
// (2, 10, 'neigh_op_top_4')
// (2, 11, 'lutff_4/out')
// (2, 11, 'sp4_h_r_8')
// (2, 12, 'neigh_op_bot_4')
// (3, 10, 'neigh_op_tnl_4')
// (3, 11, 'neigh_op_lft_4')
// (3, 11, 'sp4_h_r_21')
// (3, 12, 'neigh_op_bnl_4')
// (4, 11, 'sp4_h_r_32')
// (5, 11, 'local_g3_5')
// (5, 11, 'lutff_0/in_0')
// (5, 11, 'lutff_7/in_1')
// (5, 11, 'sp4_h_r_45')
// (6, 11, 'sp4_h_l_45')

reg n86 = 0;
// (1, 11, 'sp12_h_r_1')
// (2, 11, 'sp12_h_r_2')
// (3, 11, 'sp12_h_r_5')
// (4, 11, 'sp12_h_r_6')
// (5, 11, 'sp12_h_r_9')
// (6, 11, 'sp12_h_r_10')
// (7, 11, 'sp12_h_r_13')
// (8, 11, 'sp12_h_r_14')
// (9, 11, 'local_g0_1')
// (9, 11, 'lutff_5/in_0')
// (9, 11, 'sp12_h_r_17')
// (10, 11, 'sp12_h_r_18')
// (11, 10, 'neigh_op_tnr_7')
// (11, 11, 'neigh_op_rgt_7')
// (11, 11, 'sp12_h_r_21')
// (11, 12, 'neigh_op_bnr_7')
// (12, 10, 'neigh_op_top_7')
// (12, 11, 'lutff_7/out')
// (12, 11, 'sp12_h_r_22')
// (12, 12, 'neigh_op_bot_7')
// (13, 10, 'logic_op_tnl_7')
// (13, 11, 'logic_op_lft_7')
// (13, 11, 'span12_horz_22')
// (13, 12, 'logic_op_bnl_7')

reg n87 = 0;
// (1, 12, 'sp12_h_r_0')
// (2, 12, 'sp12_h_r_3')
// (3, 12, 'sp12_h_r_4')
// (4, 12, 'sp12_h_r_7')
// (5, 12, 'sp12_h_r_8')
// (6, 12, 'sp12_h_r_11')
// (7, 12, 'sp12_h_r_12')
// (8, 12, 'sp12_h_r_15')
// (9, 12, 'local_g0_0')
// (9, 12, 'lutff_4/in_2')
// (9, 12, 'lutff_7/in_1')
// (9, 12, 'sp12_h_r_16')
// (10, 11, 'neigh_op_tnr_6')
// (10, 12, 'neigh_op_rgt_6')
// (10, 12, 'sp12_h_r_19')
// (10, 13, 'neigh_op_bnr_6')
// (11, 11, 'neigh_op_top_6')
// (11, 12, 'lutff_6/out')
// (11, 12, 'sp12_h_r_20')
// (11, 13, 'neigh_op_bot_6')
// (12, 11, 'neigh_op_tnl_6')
// (12, 12, 'neigh_op_lft_6')
// (12, 12, 'sp12_h_r_23')
// (12, 13, 'neigh_op_bnl_6')
// (13, 12, 'span12_horz_23')

wire n88;
// (2, 3, 'sp4_h_r_8')
// (3, 2, 'neigh_op_tnr_0')
// (3, 3, 'neigh_op_rgt_0')
// (3, 3, 'sp4_h_r_21')
// (3, 4, 'neigh_op_bnr_0')
// (4, 0, 'span12_vert_20')
// (4, 1, 'sp12_v_b_20')
// (4, 2, 'neigh_op_top_0')
// (4, 2, 'sp12_v_b_19')
// (4, 2, 'sp4_r_v_b_44')
// (4, 3, 'lutff_0/out')
// (4, 3, 'sp12_v_b_16')
// (4, 3, 'sp4_h_r_32')
// (4, 3, 'sp4_r_v_b_33')
// (4, 4, 'neigh_op_bot_0')
// (4, 4, 'sp12_v_b_15')
// (4, 4, 'sp4_r_v_b_20')
// (4, 5, 'sp12_v_b_12')
// (4, 5, 'sp4_r_v_b_9')
// (4, 6, 'sp12_v_b_11')
// (4, 6, 'sp4_r_v_b_37')
// (4, 7, 'local_g2_0')
// (4, 7, 'lutff_4/in_0')
// (4, 7, 'sp12_v_b_8')
// (4, 7, 'sp4_r_v_b_24')
// (4, 8, 'sp12_v_b_7')
// (4, 8, 'sp4_r_v_b_13')
// (4, 9, 'sp12_v_b_4')
// (4, 9, 'sp4_r_v_b_0')
// (4, 10, 'local_g3_3')
// (4, 10, 'lutff_7/in_1')
// (4, 10, 'sp12_v_b_3')
// (4, 11, 'sp12_h_r_0')
// (4, 11, 'sp12_v_b_0')
// (5, 1, 'sp4_r_v_b_32')
// (5, 1, 'sp4_v_t_44')
// (5, 2, 'neigh_op_tnl_0')
// (5, 2, 'sp4_r_v_b_21')
// (5, 2, 'sp4_v_b_44')
// (5, 3, 'neigh_op_lft_0')
// (5, 3, 'sp4_h_r_45')
// (5, 3, 'sp4_r_v_b_8')
// (5, 3, 'sp4_v_b_33')
// (5, 4, 'neigh_op_bnl_0')
// (5, 4, 'sp4_v_b_20')
// (5, 5, 'sp4_v_b_9')
// (5, 5, 'sp4_v_t_37')
// (5, 6, 'sp4_v_b_37')
// (5, 7, 'sp4_v_b_24')
// (5, 8, 'local_g0_5')
// (5, 8, 'lutff_6/in_1')
// (5, 8, 'sp4_v_b_13')
// (5, 9, 'sp4_h_r_0')
// (5, 9, 'sp4_v_b_0')
// (5, 11, 'sp12_h_r_3')
// (6, 0, 'span4_vert_32')
// (6, 1, 'sp4_v_b_32')
// (6, 2, 'local_g0_5')
// (6, 2, 'lutff_2/in_3')
// (6, 2, 'sp4_v_b_21')
// (6, 3, 'sp4_h_l_45')
// (6, 3, 'sp4_v_b_8')
// (6, 9, 'sp4_h_r_13')
// (6, 11, 'sp12_h_r_4')
// (7, 9, 'local_g3_0')
// (7, 9, 'lutff_2/in_1')
// (7, 9, 'sp4_h_r_24')
// (7, 11, 'sp12_h_r_7')
// (8, 6, 'sp4_r_v_b_43')
// (8, 7, 'sp4_r_v_b_30')
// (8, 8, 'sp4_r_v_b_19')
// (8, 9, 'sp4_h_r_37')
// (8, 9, 'sp4_r_v_b_6')
// (8, 11, 'sp12_h_r_8')
// (9, 5, 'sp4_h_r_6')
// (9, 5, 'sp4_v_t_43')
// (9, 6, 'sp4_v_b_43')
// (9, 7, 'sp4_v_b_30')
// (9, 8, 'local_g0_3')
// (9, 8, 'lutff_3/in_0')
// (9, 8, 'sp4_v_b_19')
// (9, 9, 'sp4_h_l_37')
// (9, 9, 'sp4_v_b_6')
// (9, 11, 'local_g1_3')
// (9, 11, 'lutff_7/in_1')
// (9, 11, 'sp12_h_r_11')
// (10, 5, 'sp4_h_r_19')
// (10, 6, 'sp4_r_v_b_37')
// (10, 7, 'sp4_r_v_b_24')
// (10, 8, 'sp4_r_v_b_13')
// (10, 9, 'sp4_r_v_b_0')
// (10, 11, 'sp12_h_r_12')
// (11, 5, 'local_g2_6')
// (11, 5, 'lutff_1/in_1')
// (11, 5, 'sp4_h_r_30')
// (11, 5, 'sp4_h_r_6')
// (11, 5, 'sp4_v_t_37')
// (11, 6, 'sp4_v_b_37')
// (11, 7, 'local_g2_0')
// (11, 7, 'lutff_7/in_1')
// (11, 7, 'sp4_v_b_24')
// (11, 8, 'sp4_v_b_13')
// (11, 9, 'sp4_v_b_0')
// (11, 11, 'sp12_h_r_15')
// (12, 5, 'sp4_h_r_19')
// (12, 5, 'sp4_h_r_43')
// (12, 11, 'sp12_h_r_16')
// (13, 5, 'span4_horz_19')
// (13, 5, 'span4_horz_43')
// (13, 11, 'span12_horz_16')

wire n89;
// (2, 5, 'lutff_1/cout')
// (2, 5, 'lutff_2/in_3')

wire n90;
// (2, 5, 'lutff_2/cout')
// (2, 5, 'lutff_3/in_3')

wire n91;
// (2, 5, 'lutff_3/cout')
// (2, 5, 'lutff_4/in_3')

wire n92;
// (2, 5, 'lutff_4/cout')
// (2, 5, 'lutff_5/in_3')

wire n93;
// (2, 5, 'lutff_5/cout')
// (2, 5, 'lutff_6/in_3')

wire n94;
// (2, 5, 'lutff_6/cout')
// (2, 5, 'lutff_7/in_3')

reg n95 = 0;
// (2, 5, 'sp12_h_r_1')
// (3, 5, 'sp12_h_r_2')
// (4, 5, 'sp12_h_r_5')
// (5, 5, 'sp12_h_r_6')
// (6, 5, 'sp12_h_r_9')
// (7, 5, 'sp12_h_r_10')
// (8, 5, 'local_g1_5')
// (8, 5, 'lutff_1/in_3')
// (8, 5, 'sp12_h_r_13')
// (9, 5, 'sp12_h_r_14')
// (10, 4, 'neigh_op_tnr_5')
// (10, 5, 'neigh_op_rgt_5')
// (10, 5, 'sp12_h_r_17')
// (10, 5, 'sp4_r_v_b_42')
// (10, 6, 'neigh_op_bnr_5')
// (10, 6, 'sp4_r_v_b_31')
// (10, 7, 'sp4_r_v_b_18')
// (10, 8, 'sp4_r_v_b_7')
// (11, 4, 'neigh_op_top_5')
// (11, 4, 'sp4_v_t_42')
// (11, 5, 'lutff_5/out')
// (11, 5, 'sp12_h_r_18')
// (11, 5, 'sp4_v_b_42')
// (11, 6, 'neigh_op_bot_5')
// (11, 6, 'sp4_v_b_31')
// (11, 7, 'sp4_v_b_18')
// (11, 8, 'local_g1_7')
// (11, 8, 'lutff_1/in_1')
// (11, 8, 'sp4_v_b_7')
// (12, 4, 'neigh_op_tnl_5')
// (12, 5, 'neigh_op_lft_5')
// (12, 5, 'sp12_h_r_21')
// (12, 6, 'neigh_op_bnl_5')
// (13, 5, 'span12_horz_21')

wire n96;
// (2, 6, 'sp12_h_r_1')
// (3, 6, 'sp12_h_r_2')
// (4, 6, 'sp12_h_r_5')
// (5, 6, 'sp12_h_r_6')
// (6, 3, 'sp4_r_v_b_39')
// (6, 4, 'sp4_r_v_b_26')
// (6, 5, 'neigh_op_tnr_1')
// (6, 5, 'sp4_r_v_b_15')
// (6, 6, 'neigh_op_rgt_1')
// (6, 6, 'sp12_h_r_9')
// (6, 6, 'sp4_r_v_b_2')
// (6, 7, 'neigh_op_bnr_1')
// (6, 7, 'sp4_r_v_b_40')
// (6, 8, 'sp4_r_v_b_29')
// (6, 9, 'sp4_r_v_b_16')
// (6, 10, 'sp4_r_v_b_5')
// (7, 2, 'sp4_v_t_39')
// (7, 3, 'sp4_v_b_39')
// (7, 4, 'sp4_v_b_26')
// (7, 5, 'neigh_op_top_1')
// (7, 5, 'sp4_v_b_15')
// (7, 6, 'lutff_1/out')
// (7, 6, 'sp12_h_r_10')
// (7, 6, 'sp4_v_b_2')
// (7, 6, 'sp4_v_t_40')
// (7, 7, 'neigh_op_bot_1')
// (7, 7, 'sp4_v_b_40')
// (7, 8, 'sp4_v_b_29')
// (7, 9, 'local_g0_0')
// (7, 9, 'lutff_2/in_2')
// (7, 9, 'sp4_v_b_16')
// (7, 10, 'sp4_h_r_11')
// (7, 10, 'sp4_v_b_5')
// (8, 5, 'neigh_op_tnl_1')
// (8, 6, 'neigh_op_lft_1')
// (8, 6, 'sp12_h_r_13')
// (8, 7, 'neigh_op_bnl_1')
// (8, 10, 'sp4_h_r_22')
// (9, 6, 'local_g1_6')
// (9, 6, 'lutff_3/in_0')
// (9, 6, 'sp12_h_r_14')
// (9, 10, 'sp4_h_r_35')
// (10, 6, 'sp12_h_r_17')
// (10, 7, 'sp4_r_v_b_40')
// (10, 8, 'sp4_r_v_b_29')
// (10, 9, 'sp4_r_v_b_16')
// (10, 10, 'sp4_h_r_46')
// (10, 10, 'sp4_r_v_b_5')
// (11, 6, 'sp12_h_r_18')
// (11, 6, 'sp4_v_t_40')
// (11, 7, 'sp4_v_b_40')
// (11, 8, 'sp4_v_b_29')
// (11, 9, 'local_g0_0')
// (11, 9, 'lutff_2/in_2')
// (11, 9, 'sp4_v_b_16')
// (11, 10, 'sp4_h_l_46')
// (11, 10, 'sp4_v_b_5')
// (12, 6, 'sp12_h_r_21')
// (13, 6, 'span12_horz_21')

wire n97;
// (2, 8, 'sp12_h_r_1')
// (3, 8, 'sp12_h_r_2')
// (4, 8, 'sp12_h_r_5')
// (5, 8, 'sp12_h_r_6')
// (6, 7, 'neigh_op_tnr_1')
// (6, 8, 'neigh_op_rgt_1')
// (6, 8, 'sp12_h_r_9')
// (6, 9, 'neigh_op_bnr_1')
// (7, 7, 'neigh_op_top_1')
// (7, 8, 'lutff_1/out')
// (7, 8, 'sp12_h_r_10')
// (7, 9, 'neigh_op_bot_1')
// (8, 7, 'neigh_op_tnl_1')
// (8, 8, 'local_g0_5')
// (8, 8, 'local_g0_6')
// (8, 8, 'lutff_3/in_2')
// (8, 8, 'lutff_7/in_1')
// (8, 8, 'neigh_op_lft_1')
// (8, 8, 'sp12_h_r_13')
// (8, 8, 'sp4_h_r_6')
// (8, 9, 'neigh_op_bnl_1')
// (9, 8, 'sp12_h_r_14')
// (9, 8, 'sp4_h_r_19')
// (10, 8, 'sp12_h_r_17')
// (10, 8, 'sp4_h_r_30')
// (11, 8, 'sp12_h_r_18')
// (11, 8, 'sp4_h_r_43')
// (12, 8, 'sp12_h_r_21')
// (12, 8, 'sp4_h_l_43')
// (13, 8, 'span12_horz_21')

reg n98 = 0;
// (2, 9, 'sp12_h_r_0')
// (3, 8, 'neigh_op_tnr_6')
// (3, 9, 'neigh_op_rgt_6')
// (3, 9, 'sp12_h_r_3')
// (3, 10, 'neigh_op_bnr_6')
// (4, 8, 'neigh_op_top_6')
// (4, 9, 'local_g1_6')
// (4, 9, 'lutff_3/in_0')
// (4, 9, 'lutff_6/out')
// (4, 9, 'sp12_h_r_4')
// (4, 10, 'neigh_op_bot_6')
// (5, 8, 'neigh_op_tnl_6')
// (5, 9, 'local_g1_6')
// (5, 9, 'lutff_7/in_0')
// (5, 9, 'neigh_op_lft_6')
// (5, 9, 'sp12_h_r_7')
// (5, 10, 'neigh_op_bnl_6')
// (6, 9, 'local_g0_0')
// (6, 9, 'local_g1_0')
// (6, 9, 'lutff_4/in_0')
// (6, 9, 'lutff_7/in_0')
// (6, 9, 'sp12_h_r_8')
// (7, 9, 'sp12_h_r_11')
// (8, 9, 'sp12_h_r_12')
// (9, 9, 'sp12_h_r_15')
// (10, 9, 'sp12_h_r_16')
// (11, 9, 'sp12_h_r_19')
// (12, 9, 'sp12_h_r_20')
// (13, 9, 'span12_horz_20')

reg n99 = 0;
// (2, 11, 'local_g0_2')
// (2, 11, 'lutff_4/in_0')
// (2, 11, 'sp4_h_r_10')
// (3, 10, 'neigh_op_tnr_1')
// (3, 11, 'neigh_op_rgt_1')
// (3, 11, 'sp4_h_r_23')
// (3, 12, 'neigh_op_bnr_1')
// (4, 10, 'neigh_op_top_1')
// (4, 11, 'lutff_1/out')
// (4, 11, 'sp4_h_r_34')
// (4, 12, 'neigh_op_bot_1')
// (5, 10, 'neigh_op_tnl_1')
// (5, 11, 'neigh_op_lft_1')
// (5, 11, 'sp4_h_r_47')
// (5, 12, 'neigh_op_bnl_1')
// (6, 11, 'sp4_h_l_47')

reg n100 = 0;
// (2, 11, 'sp12_h_r_1')
// (3, 11, 'sp12_h_r_2')
// (4, 11, 'sp12_h_r_5')
// (5, 11, 'sp12_h_r_6')
// (6, 11, 'sp12_h_r_9')
// (7, 11, 'sp12_h_r_10')
// (8, 10, 'neigh_op_tnr_3')
// (8, 11, 'neigh_op_rgt_3')
// (8, 11, 'sp12_h_r_13')
// (8, 12, 'neigh_op_bnr_3')
// (9, 10, 'neigh_op_top_3')
// (9, 11, 'lutff_3/out')
// (9, 11, 'sp12_h_r_14')
// (9, 12, 'neigh_op_bot_3')
// (10, 10, 'neigh_op_tnl_3')
// (10, 11, 'neigh_op_lft_3')
// (10, 11, 'sp12_h_r_17')
// (10, 12, 'neigh_op_bnl_3')
// (11, 11, 'local_g0_2')
// (11, 11, 'local_g1_2')
// (11, 11, 'lutff_2/in_1')
// (11, 11, 'lutff_3/in_3')
// (11, 11, 'sp12_h_r_18')
// (12, 11, 'sp12_h_r_21')
// (13, 11, 'span12_horz_21')

reg n101 = 0;
// (2, 11, 'sp4_h_r_1')
// (3, 11, 'sp4_h_r_12')
// (4, 11, 'sp4_h_r_25')
// (5, 4, 'local_g3_0')
// (5, 4, 'lutff_5/in_0')
// (5, 4, 'sp4_r_v_b_40')
// (5, 5, 'sp4_r_v_b_29')
// (5, 6, 'sp4_r_v_b_16')
// (5, 7, 'sp4_r_v_b_5')
// (5, 8, 'sp4_r_v_b_45')
// (5, 9, 'sp4_r_v_b_32')
// (5, 10, 'sp4_r_v_b_21')
// (5, 11, 'sp4_h_r_36')
// (5, 11, 'sp4_r_v_b_8')
// (5, 12, 'local_g3_1')
// (5, 12, 'lutff_2/in_2')
// (5, 12, 'sp4_r_v_b_36')
// (5, 12, 'sp4_r_v_b_41')
// (5, 13, 'sp4_r_v_b_25')
// (5, 13, 'sp4_r_v_b_28')
// (5, 14, 'sp4_r_v_b_12')
// (5, 14, 'sp4_r_v_b_17')
// (5, 15, 'sp4_r_v_b_1')
// (5, 15, 'sp4_r_v_b_4')
// (6, 3, 'sp4_h_r_11')
// (6, 3, 'sp4_v_t_40')
// (6, 4, 'sp4_v_b_40')
// (6, 5, 'sp4_v_b_29')
// (6, 6, 'sp4_v_b_16')
// (6, 7, 'sp4_v_b_5')
// (6, 7, 'sp4_v_t_45')
// (6, 8, 'sp4_v_b_45')
// (6, 9, 'sp4_v_b_32')
// (6, 10, 'local_g0_5')
// (6, 10, 'lutff_7/in_0')
// (6, 10, 'sp4_v_b_21')
// (6, 11, 'sp4_h_l_36')
// (6, 11, 'sp4_v_b_8')
// (6, 11, 'sp4_v_t_36')
// (6, 11, 'sp4_v_t_41')
// (6, 12, 'local_g2_4')
// (6, 12, 'lutff_4/in_2')
// (6, 12, 'sp4_v_b_36')
// (6, 12, 'sp4_v_b_41')
// (6, 13, 'sp4_v_b_25')
// (6, 13, 'sp4_v_b_28')
// (6, 14, 'sp4_v_b_12')
// (6, 14, 'sp4_v_b_17')
// (6, 15, 'sp4_v_b_1')
// (6, 15, 'sp4_v_b_4')
// (7, 3, 'sp4_h_r_22')
// (8, 2, 'neigh_op_tnr_7')
// (8, 3, 'neigh_op_rgt_7')
// (8, 3, 'sp4_h_r_35')
// (8, 4, 'neigh_op_bnr_7')
// (9, 2, 'neigh_op_top_7')
// (9, 3, 'lutff_7/out')
// (9, 3, 'sp4_h_r_46')
// (9, 4, 'neigh_op_bot_7')
// (10, 2, 'neigh_op_tnl_7')
// (10, 3, 'neigh_op_lft_7')
// (10, 3, 'sp4_h_l_46')
// (10, 4, 'neigh_op_bnl_7')

wire \d_out[5] ;
// (3, 0, 'span4_horz_r_0')
// (4, 0, 'span4_horz_r_4')
// (5, 0, 'io_0/D_OUT_0')
// (5, 0, 'io_0/PAD')
// (5, 0, 'local_g0_0')
// (5, 0, 'span4_horz_r_8')
// (6, 0, 'span4_horz_r_12')
// (7, 0, 'span4_horz_l_12')
// (7, 0, 'span4_horz_r_0')
// (8, 0, 'span4_horz_r_4')
// (9, 0, 'span4_horz_r_8')
// (10, 0, 'span4_horz_r_12')
// (10, 1, 'sp4_r_v_b_25')
// (10, 2, 'sp4_r_v_b_12')
// (10, 3, 'sp4_r_v_b_1')
// (10, 4, 'sp4_r_v_b_40')
// (10, 5, 'neigh_op_tnr_0')
// (10, 5, 'sp4_r_v_b_29')
// (10, 6, 'neigh_op_rgt_0')
// (10, 6, 'sp4_r_v_b_16')
// (10, 7, 'neigh_op_bnr_0')
// (10, 7, 'sp4_r_v_b_5')
// (11, 0, 'span4_horz_l_12')
// (11, 0, 'span4_vert_25')
// (11, 1, 'sp4_v_b_25')
// (11, 2, 'sp4_v_b_12')
// (11, 3, 'sp4_v_b_1')
// (11, 3, 'sp4_v_t_40')
// (11, 4, 'sp4_v_b_40')
// (11, 5, 'neigh_op_top_0')
// (11, 5, 'sp4_v_b_29')
// (11, 6, 'lutff_0/out')
// (11, 6, 'sp4_v_b_16')
// (11, 7, 'neigh_op_bot_0')
// (11, 7, 'sp4_v_b_5')
// (12, 5, 'neigh_op_tnl_0')
// (12, 6, 'neigh_op_lft_0')
// (12, 7, 'neigh_op_bnl_0')

wire n103;
// (3, 1, 'neigh_op_tnr_5')
// (3, 2, 'neigh_op_rgt_5')
// (3, 3, 'neigh_op_bnr_5')
// (4, 1, 'neigh_op_top_5')
// (4, 2, 'local_g0_5')
// (4, 2, 'lutff_5/out')
// (4, 2, 'lutff_7/in_2')
// (4, 3, 'neigh_op_bot_5')
// (5, 1, 'neigh_op_tnl_5')
// (5, 2, 'neigh_op_lft_5')
// (5, 3, 'neigh_op_bnl_5')

wire \d_out[7] ;
// (3, 1, 'sp4_r_v_b_16')
// (3, 2, 'sp4_r_v_b_5')
// (3, 3, 'sp4_r_v_b_39')
// (3, 4, 'sp4_r_v_b_26')
// (3, 5, 'sp4_r_v_b_15')
// (3, 6, 'sp4_r_v_b_2')
// (4, 0, 'io_0/D_OUT_0')
// (4, 0, 'io_0/PAD')
// (4, 0, 'local_g0_0')
// (4, 0, 'span4_vert_16')
// (4, 1, 'sp4_v_b_16')
// (4, 2, 'sp4_v_b_5')
// (4, 2, 'sp4_v_t_39')
// (4, 3, 'sp4_v_b_39')
// (4, 4, 'sp4_v_b_26')
// (4, 5, 'neigh_op_tnr_2')
// (4, 5, 'sp4_v_b_15')
// (4, 6, 'neigh_op_rgt_2')
// (4, 6, 'sp4_h_r_9')
// (4, 6, 'sp4_v_b_2')
// (4, 7, 'neigh_op_bnr_2')
// (5, 5, 'neigh_op_top_2')
// (5, 6, 'lutff_2/out')
// (5, 6, 'sp4_h_r_20')
// (5, 7, 'neigh_op_bot_2')
// (6, 5, 'neigh_op_tnl_2')
// (6, 6, 'neigh_op_lft_2')
// (6, 6, 'sp4_h_r_33')
// (6, 7, 'neigh_op_bnl_2')
// (7, 6, 'sp4_h_r_44')
// (8, 6, 'sp4_h_l_44')

reg n105 = 0;
// (3, 3, 'neigh_op_tnr_0')
// (3, 4, 'neigh_op_rgt_0')
// (3, 5, 'neigh_op_bnr_0')
// (4, 3, 'neigh_op_top_0')
// (4, 4, 'local_g0_0')
// (4, 4, 'lutff_0/out')
// (4, 4, 'lutff_4/in_0')
// (4, 5, 'neigh_op_bot_0')
// (5, 3, 'neigh_op_tnl_0')
// (5, 4, 'neigh_op_lft_0')
// (5, 5, 'neigh_op_bnl_0')

reg n106 = 0;
// (3, 3, 'neigh_op_tnr_4')
// (3, 4, 'neigh_op_rgt_4')
// (3, 5, 'neigh_op_bnr_4')
// (4, 3, 'neigh_op_top_4')
// (4, 4, 'local_g1_4')
// (4, 4, 'lutff_4/out')
// (4, 4, 'lutff_5/in_0')
// (4, 5, 'neigh_op_bot_4')
// (5, 3, 'neigh_op_tnl_4')
// (5, 4, 'local_g1_4')
// (5, 4, 'lutff_4/in_3')
// (5, 4, 'neigh_op_lft_4')
// (5, 5, 'neigh_op_bnl_4')

reg n107 = 0;
// (3, 3, 'neigh_op_tnr_5')
// (3, 4, 'neigh_op_rgt_5')
// (3, 5, 'neigh_op_bnr_5')
// (3, 7, 'sp4_r_v_b_36')
// (3, 8, 'sp4_r_v_b_25')
// (3, 9, 'sp4_r_v_b_12')
// (3, 10, 'sp4_r_v_b_1')
// (4, 0, 'span12_vert_17')
// (4, 1, 'sp12_v_b_17')
// (4, 2, 'sp12_v_b_14')
// (4, 3, 'neigh_op_top_5')
// (4, 3, 'sp12_v_b_13')
// (4, 4, 'lutff_5/out')
// (4, 4, 'sp12_v_b_10')
// (4, 4, 'sp4_r_v_b_43')
// (4, 5, 'neigh_op_bot_5')
// (4, 5, 'sp12_v_b_9')
// (4, 5, 'sp4_r_v_b_30')
// (4, 6, 'sp12_v_b_6')
// (4, 6, 'sp4_h_r_1')
// (4, 6, 'sp4_r_v_b_19')
// (4, 6, 'sp4_v_t_36')
// (4, 7, 'sp12_v_b_5')
// (4, 7, 'sp4_r_v_b_6')
// (4, 7, 'sp4_v_b_36')
// (4, 8, 'sp12_v_b_2')
// (4, 8, 'sp4_r_v_b_44')
// (4, 8, 'sp4_v_b_25')
// (4, 9, 'sp12_v_b_1')
// (4, 9, 'sp4_r_v_b_33')
// (4, 9, 'sp4_v_b_12')
// (4, 10, 'local_g0_1')
// (4, 10, 'lutff_5/in_0')
// (4, 10, 'sp4_r_v_b_20')
// (4, 10, 'sp4_v_b_1')
// (4, 11, 'sp4_r_v_b_9')
// (5, 3, 'neigh_op_tnl_5')
// (5, 3, 'sp4_v_t_43')
// (5, 4, 'neigh_op_lft_5')
// (5, 4, 'sp4_v_b_43')
// (5, 5, 'neigh_op_bnl_5')
// (5, 5, 'sp4_v_b_30')
// (5, 6, 'sp4_h_r_12')
// (5, 6, 'sp4_v_b_19')
// (5, 7, 'sp4_v_b_6')
// (5, 7, 'sp4_v_t_44')
// (5, 8, 'sp4_v_b_44')
// (5, 9, 'sp4_v_b_33')
// (5, 10, 'sp4_v_b_20')
// (5, 11, 'sp4_h_r_9')
// (5, 11, 'sp4_v_b_9')
// (6, 6, 'local_g2_1')
// (6, 6, 'lutff_1/in_0')
// (6, 6, 'sp4_h_r_25')
// (6, 11, 'local_g0_4')
// (6, 11, 'lutff_0/in_2')
// (6, 11, 'lutff_4/in_2')
// (6, 11, 'sp4_h_r_20')
// (7, 6, 'sp4_h_r_36')
// (7, 11, 'sp4_h_r_33')
// (8, 6, 'sp4_h_l_36')
// (8, 11, 'sp4_h_r_44')
// (9, 11, 'sp4_h_l_44')

wire n108;
// (3, 5, 'neigh_op_tnr_0')
// (3, 6, 'neigh_op_rgt_0')
// (3, 7, 'neigh_op_bnr_0')
// (4, 5, 'neigh_op_top_0')
// (4, 6, 'lutff_0/out')
// (4, 7, 'neigh_op_bot_0')
// (5, 5, 'neigh_op_tnl_0')
// (5, 6, 'local_g0_0')
// (5, 6, 'lutff_0/in_2')
// (5, 6, 'neigh_op_lft_0')
// (5, 7, 'neigh_op_bnl_0')

wire n109;
// (3, 5, 'neigh_op_tnr_1')
// (3, 6, 'neigh_op_rgt_1')
// (3, 7, 'neigh_op_bnr_1')
// (4, 5, 'neigh_op_top_1')
// (4, 6, 'local_g1_1')
// (4, 6, 'lutff_0/in_0')
// (4, 6, 'lutff_1/out')
// (4, 6, 'lutff_4/in_2')
// (4, 7, 'neigh_op_bot_1')
// (5, 5, 'neigh_op_tnl_1')
// (5, 6, 'neigh_op_lft_1')
// (5, 7, 'neigh_op_bnl_1')

wire n110;
// (3, 5, 'neigh_op_tnr_2')
// (3, 6, 'neigh_op_rgt_2')
// (3, 7, 'neigh_op_bnr_2')
// (4, 5, 'neigh_op_top_2')
// (4, 6, 'local_g1_2')
// (4, 6, 'lutff_2/out')
// (4, 6, 'lutff_7/in_2')
// (4, 7, 'local_g1_2')
// (4, 7, 'lutff_0/in_1')
// (4, 7, 'lutff_4/in_1')
// (4, 7, 'neigh_op_bot_2')
// (5, 5, 'neigh_op_tnl_2')
// (5, 6, 'neigh_op_lft_2')
// (5, 7, 'neigh_op_bnl_2')

wire n111;
// (3, 5, 'neigh_op_tnr_4')
// (3, 6, 'neigh_op_rgt_4')
// (3, 7, 'neigh_op_bnr_4')
// (4, 5, 'neigh_op_top_4')
// (4, 6, 'local_g0_4')
// (4, 6, 'lutff_2/in_2')
// (4, 6, 'lutff_4/out')
// (4, 7, 'neigh_op_bot_4')
// (5, 5, 'neigh_op_tnl_4')
// (5, 6, 'neigh_op_lft_4')
// (5, 7, 'neigh_op_bnl_4')

wire \d_out[6] ;
// (3, 5, 'neigh_op_tnr_6')
// (3, 6, 'neigh_op_rgt_6')
// (3, 7, 'neigh_op_bnr_6')
// (4, 0, 'io_1/D_OUT_0')
// (4, 0, 'io_1/PAD')
// (4, 0, 'local_g0_7')
// (4, 0, 'span12_vert_23')
// (4, 1, 'sp12_v_b_23')
// (4, 2, 'sp12_v_b_20')
// (4, 3, 'sp12_v_b_19')
// (4, 4, 'sp12_v_b_16')
// (4, 5, 'neigh_op_top_6')
// (4, 5, 'sp12_v_b_15')
// (4, 6, 'lutff_6/out')
// (4, 6, 'sp12_v_b_12')
// (4, 7, 'neigh_op_bot_6')
// (4, 7, 'sp12_v_b_11')
// (4, 8, 'sp12_v_b_8')
// (4, 9, 'sp12_v_b_7')
// (4, 10, 'sp12_v_b_4')
// (4, 11, 'sp12_v_b_3')
// (4, 12, 'sp12_v_b_0')
// (5, 5, 'neigh_op_tnl_6')
// (5, 6, 'neigh_op_lft_6')
// (5, 7, 'neigh_op_bnl_6')

reg n113 = 0;
// (3, 5, 'neigh_op_tnr_7')
// (3, 6, 'neigh_op_rgt_7')
// (3, 7, 'neigh_op_bnr_7')
// (4, 1, 'sp12_v_t_22')
// (4, 2, 'sp12_v_b_22')
// (4, 3, 'sp12_v_b_21')
// (4, 4, 'local_g2_2')
// (4, 4, 'lutff_0/in_0')
// (4, 4, 'sp12_v_b_18')
// (4, 5, 'neigh_op_top_7')
// (4, 5, 'sp12_v_b_17')
// (4, 6, 'lutff_7/out')
// (4, 6, 'sp12_v_b_14')
// (4, 7, 'neigh_op_bot_7')
// (4, 7, 'sp12_v_b_13')
// (4, 8, 'sp12_v_b_10')
// (4, 9, 'sp12_v_b_9')
// (4, 10, 'sp12_v_b_6')
// (4, 11, 'sp12_v_b_5')
// (4, 12, 'sp12_v_b_2')
// (4, 13, 'sp12_v_b_1')
// (5, 5, 'neigh_op_tnl_7')
// (5, 6, 'neigh_op_lft_7')
// (5, 7, 'neigh_op_bnl_7')

reg n114 = 0;
// (3, 5, 'sp12_h_r_0')
// (4, 5, 'sp12_h_r_3')
// (5, 5, 'sp12_h_r_4')
// (6, 5, 'sp12_h_r_7')
// (7, 5, 'sp12_h_r_8')
// (8, 4, 'neigh_op_tnr_2')
// (8, 5, 'neigh_op_rgt_2')
// (8, 5, 'sp12_h_r_11')
// (8, 6, 'neigh_op_bnr_2')
// (9, 4, 'neigh_op_top_2')
// (9, 5, 'lutff_2/out')
// (9, 5, 'sp12_h_r_12')
// (9, 6, 'neigh_op_bot_2')
// (10, 4, 'neigh_op_tnl_2')
// (10, 5, 'neigh_op_lft_2')
// (10, 5, 'sp12_h_r_15')
// (10, 6, 'neigh_op_bnl_2')
// (11, 5, 'local_g1_0')
// (11, 5, 'lutff_5/in_0')
// (11, 5, 'sp12_h_r_16')
// (12, 5, 'sp12_h_r_19')
// (13, 5, 'span12_horz_19')

wire n115;
// (3, 5, 'sp12_h_r_1')
// (4, 5, 'sp12_h_r_2')
// (5, 5, 'sp12_h_r_5')
// (6, 5, 'sp12_h_r_6')
// (7, 4, 'neigh_op_tnr_1')
// (7, 5, 'neigh_op_rgt_1')
// (7, 5, 'sp12_h_r_9')
// (7, 5, 'sp4_h_r_4')
// (7, 6, 'neigh_op_bnr_1')
// (8, 4, 'neigh_op_top_1')
// (8, 5, 'lutff_1/out')
// (8, 5, 'sp12_h_r_10')
// (8, 5, 'sp4_h_r_17')
// (8, 6, 'neigh_op_bot_1')
// (9, 4, 'neigh_op_tnl_1')
// (9, 5, 'neigh_op_lft_1')
// (9, 5, 'sp12_h_r_13')
// (9, 5, 'sp4_h_r_28')
// (9, 6, 'neigh_op_bnl_1')
// (10, 2, 'sp4_r_v_b_41')
// (10, 3, 'sp4_r_v_b_28')
// (10, 4, 'sp4_r_v_b_17')
// (10, 5, 'sp12_h_r_14')
// (10, 5, 'sp4_h_r_41')
// (10, 5, 'sp4_r_v_b_4')
// (10, 6, 'sp4_r_v_b_42')
// (10, 7, 'sp4_r_v_b_31')
// (10, 8, 'sp4_r_v_b_18')
// (10, 9, 'sp4_r_v_b_7')
// (11, 1, 'sp4_v_t_41')
// (11, 2, 'sp4_v_b_41')
// (11, 3, 'sp4_v_b_28')
// (11, 4, 'local_g0_1')
// (11, 4, 'lutff_5/in_0')
// (11, 4, 'sp4_v_b_17')
// (11, 5, 'local_g0_1')
// (11, 5, 'lutff_1/in_2')
// (11, 5, 'sp12_h_r_17')
// (11, 5, 'sp4_h_l_41')
// (11, 5, 'sp4_v_b_4')
// (11, 5, 'sp4_v_t_42')
// (11, 6, 'sp4_v_b_42')
// (11, 7, 'sp4_v_b_31')
// (11, 8, 'local_g0_2')
// (11, 8, 'lutff_2/in_2')
// (11, 8, 'sp4_v_b_18')
// (11, 9, 'sp4_v_b_7')
// (12, 5, 'sp12_h_r_18')
// (13, 5, 'span12_horz_18')

reg n116 = 0;
// (3, 6, 'neigh_op_tnr_0')
// (3, 7, 'neigh_op_rgt_0')
// (3, 8, 'neigh_op_bnr_0')
// (4, 6, 'local_g0_0')
// (4, 6, 'lutff_6/in_2')
// (4, 6, 'neigh_op_top_0')
// (4, 7, 'lutff_0/out')
// (4, 8, 'neigh_op_bot_0')
// (5, 6, 'neigh_op_tnl_0')
// (5, 7, 'neigh_op_lft_0')
// (5, 8, 'neigh_op_bnl_0')

reg n117 = 0;
// (3, 6, 'neigh_op_tnr_1')
// (3, 7, 'neigh_op_rgt_1')
// (3, 8, 'neigh_op_bnr_1')
// (4, 6, 'neigh_op_top_1')
// (4, 7, 'local_g0_1')
// (4, 7, 'lutff_1/out')
// (4, 7, 'lutff_3/in_0')
// (4, 8, 'neigh_op_bot_1')
// (5, 6, 'neigh_op_tnl_1')
// (5, 7, 'neigh_op_lft_1')
// (5, 8, 'neigh_op_bnl_1')

reg n118 = 0;
// (3, 6, 'neigh_op_tnr_2')
// (3, 7, 'neigh_op_rgt_2')
// (3, 8, 'neigh_op_bnr_2')
// (4, 6, 'neigh_op_top_2')
// (4, 7, 'local_g3_2')
// (4, 7, 'lutff_1/in_0')
// (4, 7, 'lutff_2/out')
// (4, 8, 'neigh_op_bot_2')
// (5, 6, 'neigh_op_tnl_2')
// (5, 7, 'neigh_op_lft_2')
// (5, 8, 'neigh_op_bnl_2')

reg n119 = 0;
// (3, 6, 'neigh_op_tnr_3')
// (3, 7, 'neigh_op_rgt_3')
// (3, 8, 'neigh_op_bnr_3')
// (4, 5, 'sp4_r_v_b_47')
// (4, 6, 'local_g0_1')
// (4, 6, 'local_g1_3')
// (4, 6, 'lutff_6/in_1')
// (4, 6, 'lutff_7/in_3')
// (4, 6, 'neigh_op_top_3')
// (4, 6, 'sp4_r_v_b_34')
// (4, 7, 'local_g0_3')
// (4, 7, 'local_g1_3')
// (4, 7, 'lutff_0/in_3')
// (4, 7, 'lutff_3/out')
// (4, 7, 'lutff_4/in_2')
// (4, 7, 'sp4_r_v_b_23')
// (4, 8, 'neigh_op_bot_3')
// (4, 8, 'sp4_r_v_b_10')
// (5, 4, 'sp4_v_t_47')
// (5, 5, 'sp4_v_b_47')
// (5, 6, 'neigh_op_tnl_3')
// (5, 6, 'sp4_v_b_34')
// (5, 7, 'neigh_op_lft_3')
// (5, 7, 'sp4_v_b_23')
// (5, 8, 'neigh_op_bnl_3')
// (5, 8, 'sp4_v_b_10')

reg n120 = 0;
// (3, 6, 'neigh_op_tnr_4')
// (3, 7, 'neigh_op_rgt_4')
// (3, 8, 'neigh_op_bnr_4')
// (4, 6, 'neigh_op_top_4')
// (4, 7, 'local_g0_4')
// (4, 7, 'lutff_2/in_0')
// (4, 7, 'lutff_4/out')
// (4, 8, 'neigh_op_bot_4')
// (5, 6, 'neigh_op_tnl_4')
// (5, 7, 'neigh_op_lft_4')
// (5, 8, 'neigh_op_bnl_4')

reg n121 = 0;
// (3, 6, 'neigh_op_tnr_5')
// (3, 7, 'neigh_op_rgt_5')
// (3, 8, 'neigh_op_bnr_5')
// (4, 6, 'neigh_op_top_5')
// (4, 7, 'local_g0_5')
// (4, 7, 'lutff_4/in_3')
// (4, 7, 'lutff_5/out')
// (4, 8, 'neigh_op_bot_5')
// (5, 6, 'neigh_op_tnl_5')
// (5, 7, 'neigh_op_lft_5')
// (5, 8, 'neigh_op_bnl_5')

wire n122;
// (3, 6, 'sp4_h_r_2')
// (4, 6, 'sp4_h_r_15')
// (5, 6, 'sp4_h_r_26')
// (6, 6, 'sp4_h_r_39')
// (6, 7, 'sp4_r_v_b_39')
// (6, 7, 'sp4_r_v_b_45')
// (6, 8, 'local_g0_2')
// (6, 8, 'local_g0_3')
// (6, 8, 'lutff_3/in_3')
// (6, 8, 'lutff_4/in_2')
// (6, 8, 'lutff_6/in_3')
// (6, 8, 'sp4_r_v_b_26')
// (6, 8, 'sp4_r_v_b_32')
// (6, 9, 'local_g2_4')
// (6, 9, 'lutff_0/in_2')
// (6, 9, 'neigh_op_tnr_4')
// (6, 9, 'sp4_r_v_b_15')
// (6, 9, 'sp4_r_v_b_21')
// (6, 10, 'neigh_op_rgt_4')
// (6, 10, 'sp4_r_v_b_2')
// (6, 10, 'sp4_r_v_b_8')
// (6, 11, 'neigh_op_bnr_4')
// (7, 6, 'sp4_h_l_39')
// (7, 6, 'sp4_v_t_39')
// (7, 6, 'sp4_v_t_45')
// (7, 7, 'sp4_v_b_39')
// (7, 7, 'sp4_v_b_45')
// (7, 8, 'sp4_v_b_26')
// (7, 8, 'sp4_v_b_32')
// (7, 9, 'neigh_op_top_4')
// (7, 9, 'sp4_v_b_15')
// (7, 9, 'sp4_v_b_21')
// (7, 10, 'lutff_4/out')
// (7, 10, 'sp4_v_b_2')
// (7, 10, 'sp4_v_b_8')
// (7, 11, 'neigh_op_bot_4')
// (8, 9, 'neigh_op_tnl_4')
// (8, 10, 'neigh_op_lft_4')
// (8, 11, 'neigh_op_bnl_4')

reg n123 = 0;
// (3, 7, 'neigh_op_tnr_1')
// (3, 8, 'neigh_op_rgt_1')
// (3, 9, 'neigh_op_bnr_1')
// (4, 7, 'neigh_op_top_1')
// (4, 8, 'local_g0_1')
// (4, 8, 'lutff_1/out')
// (4, 8, 'lutff_5/in_0')
// (4, 9, 'neigh_op_bot_1')
// (5, 7, 'neigh_op_tnl_1')
// (5, 8, 'neigh_op_lft_1')
// (5, 9, 'neigh_op_bnl_1')

reg n124 = 0;
// (3, 7, 'neigh_op_tnr_2')
// (3, 8, 'neigh_op_rgt_2')
// (3, 9, 'neigh_op_bnr_2')
// (4, 7, 'neigh_op_top_2')
// (4, 8, 'lutff_2/out')
// (4, 8, 'sp4_h_r_4')
// (4, 9, 'neigh_op_bot_2')
// (5, 7, 'neigh_op_tnl_2')
// (5, 8, 'local_g0_1')
// (5, 8, 'lutff_7/in_0')
// (5, 8, 'neigh_op_lft_2')
// (5, 8, 'sp4_h_r_17')
// (5, 9, 'neigh_op_bnl_2')
// (6, 8, 'sp4_h_r_28')
// (7, 8, 'sp4_h_r_41')
// (8, 8, 'sp4_h_l_41')

reg n125 = 0;
// (3, 7, 'neigh_op_tnr_4')
// (3, 8, 'neigh_op_rgt_4')
// (3, 9, 'neigh_op_bnr_4')
// (4, 7, 'local_g1_4')
// (4, 7, 'lutff_5/in_0')
// (4, 7, 'neigh_op_top_4')
// (4, 8, 'lutff_4/out')
// (4, 9, 'neigh_op_bot_4')
// (5, 7, 'neigh_op_tnl_4')
// (5, 8, 'neigh_op_lft_4')
// (5, 9, 'neigh_op_bnl_4')

reg n126 = 0;
// (3, 7, 'neigh_op_tnr_5')
// (3, 8, 'neigh_op_rgt_5')
// (3, 9, 'neigh_op_bnr_5')
// (4, 7, 'neigh_op_top_5')
// (4, 8, 'local_g1_5')
// (4, 8, 'lutff_4/in_0')
// (4, 8, 'lutff_5/out')
// (4, 9, 'neigh_op_bot_5')
// (5, 7, 'neigh_op_tnl_5')
// (5, 8, 'neigh_op_lft_5')
// (5, 9, 'neigh_op_bnl_5')

reg n127 = 0;
// (3, 8, 'neigh_op_tnr_0')
// (3, 9, 'neigh_op_rgt_0')
// (3, 10, 'neigh_op_bnr_0')
// (4, 8, 'neigh_op_top_0')
// (4, 9, 'local_g1_0')
// (4, 9, 'lutff_0/out')
// (4, 9, 'lutff_7/in_0')
// (4, 10, 'neigh_op_bot_0')
// (5, 8, 'neigh_op_tnl_0')
// (5, 9, 'neigh_op_lft_0')
// (5, 10, 'neigh_op_bnl_0')

reg n128 = 0;
// (3, 8, 'neigh_op_tnr_4')
// (3, 9, 'neigh_op_rgt_4')
// (3, 10, 'neigh_op_bnr_4')
// (4, 8, 'neigh_op_top_4')
// (4, 9, 'local_g2_4')
// (4, 9, 'lutff_4/out')
// (4, 9, 'lutff_6/in_0')
// (4, 10, 'neigh_op_bot_4')
// (5, 8, 'neigh_op_tnl_4')
// (5, 9, 'neigh_op_lft_4')
// (5, 10, 'neigh_op_bnl_4')

reg n129 = 0;
// (3, 8, 'neigh_op_tnr_5')
// (3, 9, 'neigh_op_rgt_5')
// (3, 10, 'neigh_op_bnr_5')
// (4, 8, 'neigh_op_top_5')
// (4, 9, 'local_g1_5')
// (4, 9, 'lutff_0/in_0')
// (4, 9, 'lutff_5/out')
// (4, 10, 'neigh_op_bot_5')
// (5, 8, 'neigh_op_tnl_5')
// (5, 9, 'neigh_op_lft_5')
// (5, 10, 'neigh_op_bnl_5')

reg n130 = 0;
// (3, 9, 'neigh_op_tnr_0')
// (3, 10, 'neigh_op_rgt_0')
// (3, 11, 'neigh_op_bnr_0')
// (4, 9, 'neigh_op_top_0')
// (4, 10, 'local_g2_0')
// (4, 10, 'lutff_0/out')
// (4, 10, 'lutff_7/in_3')
// (4, 11, 'neigh_op_bot_0')
// (5, 9, 'neigh_op_tnl_0')
// (5, 10, 'neigh_op_lft_0')
// (5, 11, 'neigh_op_bnl_0')

reg n131 = 0;
// (3, 9, 'neigh_op_tnr_1')
// (3, 10, 'neigh_op_rgt_1')
// (3, 11, 'neigh_op_bnr_1')
// (4, 7, 'sp4_r_v_b_38')
// (4, 8, 'local_g0_3')
// (4, 8, 'lutff_1/in_0')
// (4, 8, 'sp4_r_v_b_27')
// (4, 9, 'neigh_op_top_1')
// (4, 9, 'sp4_r_v_b_14')
// (4, 10, 'lutff_1/out')
// (4, 10, 'sp4_r_v_b_3')
// (4, 11, 'neigh_op_bot_1')
// (5, 6, 'sp4_v_t_38')
// (5, 7, 'sp4_v_b_38')
// (5, 8, 'sp4_v_b_27')
// (5, 9, 'neigh_op_tnl_1')
// (5, 9, 'sp4_v_b_14')
// (5, 10, 'neigh_op_lft_1')
// (5, 10, 'sp4_v_b_3')
// (5, 11, 'neigh_op_bnl_1')

reg n132 = 0;
// (3, 9, 'neigh_op_tnr_2')
// (3, 10, 'neigh_op_rgt_2')
// (3, 11, 'neigh_op_bnr_2')
// (4, 9, 'neigh_op_top_2')
// (4, 10, 'lutff_2/out')
// (4, 11, 'neigh_op_bot_2')
// (5, 9, 'neigh_op_tnl_2')
// (5, 10, 'local_g0_2')
// (5, 10, 'lutff_4/in_0')
// (5, 10, 'neigh_op_lft_2')
// (5, 11, 'neigh_op_bnl_2')

reg n133 = 0;
// (3, 9, 'neigh_op_tnr_4')
// (3, 10, 'neigh_op_rgt_4')
// (3, 11, 'neigh_op_bnr_4')
// (4, 9, 'neigh_op_top_4')
// (4, 10, 'local_g0_4')
// (4, 10, 'lutff_4/out')
// (4, 10, 'lutff_6/in_0')
// (4, 11, 'neigh_op_bot_4')
// (5, 9, 'neigh_op_tnl_4')
// (5, 10, 'neigh_op_lft_4')
// (5, 11, 'neigh_op_bnl_4')

reg n134 = 0;
// (3, 9, 'neigh_op_tnr_5')
// (3, 10, 'neigh_op_rgt_5')
// (3, 11, 'neigh_op_bnr_5')
// (4, 9, 'neigh_op_top_5')
// (4, 10, 'local_g1_5')
// (4, 10, 'lutff_4/in_0')
// (4, 10, 'lutff_5/out')
// (4, 11, 'neigh_op_bot_5')
// (5, 9, 'neigh_op_tnl_5')
// (5, 10, 'neigh_op_lft_5')
// (5, 11, 'neigh_op_bnl_5')

reg n135 = 0;
// (3, 9, 'neigh_op_tnr_6')
// (3, 10, 'neigh_op_rgt_6')
// (3, 11, 'neigh_op_bnr_6')
// (4, 9, 'neigh_op_top_6')
// (4, 10, 'local_g1_6')
// (4, 10, 'lutff_1/in_0')
// (4, 10, 'lutff_6/out')
// (4, 11, 'neigh_op_bot_6')
// (5, 9, 'neigh_op_tnl_6')
// (5, 10, 'neigh_op_lft_6')
// (5, 11, 'neigh_op_bnl_6')

reg n136 = 0;
// (3, 9, 'neigh_op_tnr_7')
// (3, 10, 'neigh_op_rgt_7')
// (3, 11, 'neigh_op_bnr_7')
// (4, 9, 'neigh_op_top_7')
// (4, 10, 'local_g1_7')
// (4, 10, 'lutff_2/in_0')
// (4, 10, 'lutff_7/out')
// (4, 11, 'neigh_op_bot_7')
// (5, 9, 'neigh_op_tnl_7')
// (5, 10, 'neigh_op_lft_7')
// (5, 11, 'neigh_op_bnl_7')

wire n137;
// (3, 9, 'sp12_h_r_1')
// (4, 9, 'sp12_h_r_2')
// (5, 9, 'sp12_h_r_5')
// (6, 9, 'sp12_h_r_6')
// (7, 8, 'neigh_op_tnr_1')
// (7, 9, 'neigh_op_rgt_1')
// (7, 9, 'sp12_h_r_9')
// (7, 10, 'neigh_op_bnr_1')
// (8, 8, 'neigh_op_top_1')
// (8, 9, 'lutff_1/out')
// (8, 9, 'sp12_h_r_10')
// (8, 10, 'neigh_op_bot_1')
// (9, 8, 'neigh_op_tnl_1')
// (9, 9, 'neigh_op_lft_1')
// (9, 9, 'sp12_h_r_13')
// (9, 10, 'neigh_op_bnl_1')
// (10, 9, 'sp12_h_r_14')
// (11, 9, 'local_g1_1')
// (11, 9, 'lutff_1/in_3')
// (11, 9, 'lutff_4/in_2')
// (11, 9, 'sp12_h_r_17')
// (12, 9, 'sp12_h_r_18')
// (13, 9, 'span12_horz_18')

reg n138 = 0;
// (3, 10, 'neigh_op_tnr_0')
// (3, 11, 'neigh_op_rgt_0')
// (3, 12, 'neigh_op_bnr_0')
// (4, 10, 'neigh_op_top_0')
// (4, 11, 'local_g1_0')
// (4, 11, 'lutff_0/out')
// (4, 11, 'lutff_3/in_0')
// (4, 12, 'neigh_op_bot_0')
// (5, 10, 'neigh_op_tnl_0')
// (5, 11, 'neigh_op_lft_0')
// (5, 12, 'neigh_op_bnl_0')

reg n139 = 0;
// (3, 10, 'neigh_op_tnr_2')
// (3, 11, 'neigh_op_rgt_2')
// (3, 12, 'neigh_op_bnr_2')
// (4, 10, 'neigh_op_top_2')
// (4, 11, 'local_g1_2')
// (4, 11, 'lutff_1/in_0')
// (4, 11, 'lutff_2/out')
// (4, 12, 'neigh_op_bot_2')
// (5, 10, 'neigh_op_tnl_2')
// (5, 11, 'neigh_op_lft_2')
// (5, 12, 'neigh_op_bnl_2')

reg n140 = 0;
// (3, 10, 'neigh_op_tnr_3')
// (3, 11, 'neigh_op_rgt_3')
// (3, 12, 'neigh_op_bnr_3')
// (4, 10, 'local_g1_3')
// (4, 10, 'lutff_0/in_0')
// (4, 10, 'neigh_op_top_3')
// (4, 11, 'lutff_3/out')
// (4, 12, 'neigh_op_bot_3')
// (5, 10, 'neigh_op_tnl_3')
// (5, 11, 'neigh_op_lft_3')
// (5, 12, 'neigh_op_bnl_3')

reg n141 = 0;
// (3, 10, 'neigh_op_tnr_7')
// (3, 11, 'neigh_op_rgt_7')
// (3, 12, 'neigh_op_bnr_7')
// (4, 10, 'neigh_op_top_7')
// (4, 11, 'local_g1_7')
// (4, 11, 'lutff_0/in_0')
// (4, 11, 'lutff_7/out')
// (4, 12, 'neigh_op_bot_7')
// (5, 10, 'neigh_op_tnl_7')
// (5, 11, 'neigh_op_lft_7')
// (5, 12, 'neigh_op_bnl_7')

reg n142 = 0;
// (3, 11, 'neigh_op_tnr_0')
// (3, 12, 'neigh_op_rgt_0')
// (3, 13, 'neigh_op_bnr_0')
// (4, 11, 'local_g0_0')
// (4, 11, 'lutff_4/in_0')
// (4, 11, 'neigh_op_top_0')
// (4, 12, 'lutff_0/out')
// (4, 13, 'neigh_op_bot_0')
// (5, 11, 'neigh_op_tnl_0')
// (5, 12, 'neigh_op_lft_0')
// (5, 13, 'neigh_op_bnl_0')

reg n143 = 0;
// (3, 11, 'neigh_op_tnr_1')
// (3, 12, 'neigh_op_rgt_1')
// (3, 13, 'neigh_op_bnr_1')
// (4, 11, 'neigh_op_top_1')
// (4, 12, 'local_g1_1')
// (4, 12, 'lutff_1/out')
// (4, 12, 'lutff_6/in_0')
// (4, 13, 'neigh_op_bot_1')
// (5, 11, 'neigh_op_tnl_1')
// (5, 12, 'neigh_op_lft_1')
// (5, 13, 'neigh_op_bnl_1')

reg n144 = 0;
// (3, 11, 'neigh_op_tnr_2')
// (3, 12, 'neigh_op_rgt_2')
// (3, 13, 'neigh_op_bnr_2')
// (4, 11, 'neigh_op_top_2')
// (4, 12, 'local_g0_2')
// (4, 12, 'lutff_0/in_0')
// (4, 12, 'lutff_2/out')
// (4, 13, 'neigh_op_bot_2')
// (5, 11, 'neigh_op_tnl_2')
// (5, 12, 'neigh_op_lft_2')
// (5, 13, 'neigh_op_bnl_2')

reg n145 = 0;
// (3, 11, 'neigh_op_tnr_6')
// (3, 12, 'neigh_op_rgt_6')
// (3, 13, 'neigh_op_bnr_6')
// (4, 11, 'local_g1_6')
// (4, 11, 'lutff_7/in_0')
// (4, 11, 'neigh_op_top_6')
// (4, 12, 'lutff_6/out')
// (4, 13, 'neigh_op_bot_6')
// (5, 11, 'neigh_op_tnl_6')
// (5, 12, 'neigh_op_lft_6')
// (5, 13, 'neigh_op_bnl_6')

reg n146 = 0;
// (3, 11, 'sp12_h_r_0')
// (4, 11, 'sp12_h_r_3')
// (5, 11, 'sp12_h_r_4')
// (6, 11, 'sp12_h_r_7')
// (7, 11, 'sp12_h_r_8')
// (8, 11, 'local_g0_3')
// (8, 11, 'lutff_6/in_1')
// (8, 11, 'sp12_h_r_11')
// (9, 11, 'sp12_h_r_12')
// (10, 10, 'neigh_op_tnr_4')
// (10, 11, 'neigh_op_rgt_4')
// (10, 11, 'sp12_h_r_15')
// (10, 12, 'neigh_op_bnr_4')
// (11, 10, 'neigh_op_top_4')
// (11, 11, 'lutff_4/out')
// (11, 11, 'sp12_h_r_16')
// (11, 12, 'neigh_op_bot_4')
// (12, 10, 'neigh_op_tnl_4')
// (12, 11, 'neigh_op_lft_4')
// (12, 11, 'sp12_h_r_19')
// (12, 12, 'neigh_op_bnl_4')
// (13, 11, 'span12_horz_19')

wire n147;
// (3, 12, 'sp12_h_r_1')
// (4, 12, 'sp12_h_r_2')
// (5, 12, 'local_g0_5')
// (5, 12, 'lutff_2/in_1')
// (5, 12, 'sp12_h_r_5')
// (6, 12, 'local_g1_6')
// (6, 12, 'lutff_4/in_1')
// (6, 12, 'sp12_h_r_6')
// (7, 11, 'neigh_op_tnr_1')
// (7, 12, 'neigh_op_rgt_1')
// (7, 12, 'sp12_h_r_9')
// (7, 13, 'neigh_op_bnr_1')
// (8, 11, 'neigh_op_top_1')
// (8, 12, 'lutff_1/out')
// (8, 12, 'sp12_h_r_10')
// (8, 13, 'neigh_op_bot_1')
// (9, 11, 'neigh_op_tnl_1')
// (9, 12, 'neigh_op_lft_1')
// (9, 12, 'sp12_h_r_13')
// (9, 13, 'neigh_op_bnl_1')
// (10, 12, 'sp12_h_r_14')
// (11, 12, 'sp12_h_r_17')
// (12, 12, 'sp12_h_r_18')
// (13, 12, 'span12_horz_18')

reg n148 = 0;
// (4, 2, 'sp4_r_v_b_46')
// (4, 3, 'sp4_r_v_b_35')
// (4, 4, 'sp4_r_v_b_22')
// (4, 5, 'sp4_r_v_b_11')
// (4, 6, 'sp4_r_v_b_46')
// (4, 7, 'neigh_op_tnr_3')
// (4, 7, 'sp4_r_v_b_35')
// (4, 8, 'neigh_op_rgt_3')
// (4, 8, 'sp4_r_v_b_22')
// (4, 8, 'sp4_r_v_b_38')
// (4, 9, 'local_g2_3')
// (4, 9, 'lutff_5/in_0')
// (4, 9, 'neigh_op_bnr_3')
// (4, 9, 'sp4_r_v_b_11')
// (4, 9, 'sp4_r_v_b_27')
// (4, 10, 'sp4_r_v_b_14')
// (4, 11, 'sp4_r_v_b_3')
// (5, 1, 'sp4_v_t_46')
// (5, 2, 'sp4_v_b_46')
// (5, 3, 'sp4_v_b_35')
// (5, 4, 'sp4_v_b_22')
// (5, 5, 'local_g0_3')
// (5, 5, 'lutff_7/in_0')
// (5, 5, 'sp4_v_b_11')
// (5, 5, 'sp4_v_t_46')
// (5, 6, 'sp4_v_b_46')
// (5, 7, 'neigh_op_top_3')
// (5, 7, 'sp4_v_b_35')
// (5, 7, 'sp4_v_t_38')
// (5, 8, 'lutff_3/out')
// (5, 8, 'sp4_v_b_22')
// (5, 8, 'sp4_v_b_38')
// (5, 9, 'neigh_op_bot_3')
// (5, 9, 'sp4_v_b_11')
// (5, 9, 'sp4_v_b_27')
// (5, 10, 'local_g0_6')
// (5, 10, 'local_g1_6')
// (5, 10, 'lutff_2/in_2')
// (5, 10, 'lutff_7/in_2')
// (5, 10, 'sp4_v_b_14')
// (5, 11, 'sp4_v_b_3')
// (6, 7, 'neigh_op_tnl_3')
// (6, 8, 'neigh_op_lft_3')
// (6, 9, 'neigh_op_bnl_3')

wire n149;
// (4, 3, 'neigh_op_tnr_0')
// (4, 4, 'neigh_op_rgt_0')
// (4, 5, 'neigh_op_bnr_0')
// (5, 3, 'neigh_op_top_0')
// (5, 4, 'lutff_0/out')
// (5, 4, 'sp4_h_r_0')
// (5, 5, 'neigh_op_bot_0')
// (6, 3, 'local_g3_0')
// (6, 3, 'lutff_0/in_3')
// (6, 3, 'neigh_op_tnl_0')
// (6, 4, 'local_g1_0')
// (6, 4, 'local_g1_5')
// (6, 4, 'lutff_1/in_3')
// (6, 4, 'lutff_5/in_2')
// (6, 4, 'neigh_op_lft_0')
// (6, 4, 'sp4_h_r_13')
// (6, 5, 'neigh_op_bnl_0')
// (7, 4, 'sp4_h_r_24')
// (8, 4, 'sp4_h_r_37')
// (9, 4, 'sp4_h_l_37')

wire n150;
// (4, 3, 'neigh_op_tnr_4')
// (4, 4, 'neigh_op_rgt_4')
// (4, 5, 'neigh_op_bnr_4')
// (5, 3, 'neigh_op_top_4')
// (5, 4, 'lutff_4/out')
// (5, 5, 'neigh_op_bot_4')
// (6, 3, 'neigh_op_tnl_4')
// (6, 4, 'local_g1_4')
// (6, 4, 'lutff_5/in_0')
// (6, 4, 'lutff_7/in_2')
// (6, 4, 'neigh_op_lft_4')
// (6, 5, 'neigh_op_bnl_4')

reg n151 = 0;
// (4, 3, 'neigh_op_tnr_5')
// (4, 4, 'neigh_op_rgt_5')
// (4, 5, 'neigh_op_bnr_5')
// (5, 3, 'neigh_op_top_5')
// (5, 4, 'local_g0_5')
// (5, 4, 'lutff_0/in_3')
// (5, 4, 'lutff_5/out')
// (5, 5, 'neigh_op_bot_5')
// (6, 3, 'neigh_op_tnl_5')
// (6, 4, 'neigh_op_lft_5')
// (6, 5, 'neigh_op_bnl_5')

wire n152;
// (4, 3, 'sp12_h_r_0')
// (5, 2, 'neigh_op_tnr_6')
// (5, 3, 'neigh_op_rgt_6')
// (5, 3, 'sp12_h_r_3')
// (5, 4, 'neigh_op_bnr_6')
// (6, 2, 'local_g1_6')
// (6, 2, 'lutff_7/in_2')
// (6, 2, 'neigh_op_top_6')
// (6, 3, 'lutff_6/out')
// (6, 3, 'sp12_h_r_4')
// (6, 4, 'neigh_op_bot_6')
// (7, 2, 'local_g3_6')
// (7, 2, 'lutff_0/in_1')
// (7, 2, 'lutff_6/in_1')
// (7, 2, 'neigh_op_tnl_6')
// (7, 3, 'neigh_op_lft_6')
// (7, 3, 'sp12_h_r_7')
// (7, 4, 'neigh_op_bnl_6')
// (8, 3, 'local_g0_0')
// (8, 3, 'lutff_6/in_0')
// (8, 3, 'sp12_h_r_8')
// (9, 3, 'sp12_h_r_11')
// (10, 3, 'sp12_h_r_12')
// (11, 3, 'sp12_h_r_15')
// (12, 3, 'sp12_h_r_16')
// (13, 3, 'span12_horz_16')

wire n153;
// (4, 4, 'neigh_op_tnr_1')
// (4, 5, 'neigh_op_rgt_1')
// (4, 6, 'neigh_op_bnr_1')
// (5, 4, 'neigh_op_top_1')
// (5, 5, 'local_g1_1')
// (5, 5, 'lutff_1/out')
// (5, 5, 'lutff_6/in_2')
// (5, 6, 'neigh_op_bot_1')
// (6, 4, 'neigh_op_tnl_1')
// (6, 5, 'neigh_op_lft_1')
// (6, 6, 'neigh_op_bnl_1')

wire n154;
// (4, 4, 'neigh_op_tnr_2')
// (4, 5, 'neigh_op_rgt_2')
// (4, 6, 'neigh_op_bnr_2')
// (5, 4, 'neigh_op_top_2')
// (5, 5, 'local_g0_2')
// (5, 5, 'local_g1_2')
// (5, 5, 'lutff_2/out')
// (5, 5, 'lutff_3/in_3')
// (5, 5, 'lutff_6/in_3')
// (5, 6, 'neigh_op_bot_2')
// (6, 4, 'neigh_op_tnl_2')
// (6, 5, 'neigh_op_lft_2')
// (6, 6, 'neigh_op_bnl_2')

wire n155;
// (4, 4, 'neigh_op_tnr_3')
// (4, 5, 'neigh_op_rgt_3')
// (4, 6, 'neigh_op_bnr_3')
// (5, 4, 'neigh_op_top_3')
// (5, 5, 'lutff_3/out')
// (5, 5, 'sp4_r_v_b_39')
// (5, 6, 'neigh_op_bot_3')
// (5, 6, 'sp4_r_v_b_26')
// (5, 7, 'sp4_r_v_b_15')
// (5, 8, 'sp4_r_v_b_2')
// (6, 4, 'neigh_op_tnl_3')
// (6, 4, 'sp4_h_r_2')
// (6, 4, 'sp4_v_t_39')
// (6, 5, 'neigh_op_lft_3')
// (6, 5, 'sp4_v_b_39')
// (6, 6, 'neigh_op_bnl_3')
// (6, 6, 'sp4_v_b_26')
// (6, 7, 'sp4_v_b_15')
// (6, 8, 'sp4_v_b_2')
// (7, 4, 'local_g0_7')
// (7, 4, 'local_g1_7')
// (7, 4, 'lutff_0/in_2')
// (7, 4, 'lutff_2/in_3')
// (7, 4, 'lutff_3/in_1')
// (7, 4, 'lutff_6/in_2')
// (7, 4, 'sp4_h_r_15')
// (8, 4, 'sp4_h_r_26')
// (9, 4, 'sp4_h_r_39')
// (10, 4, 'sp4_h_l_39')

wire n156;
// (4, 4, 'neigh_op_tnr_4')
// (4, 5, 'neigh_op_rgt_4')
// (4, 6, 'neigh_op_bnr_4')
// (5, 4, 'neigh_op_top_4')
// (5, 5, 'local_g3_4')
// (5, 5, 'lutff_4/out')
// (5, 5, 'lutff_6/in_1')
// (5, 6, 'neigh_op_bot_4')
// (6, 4, 'neigh_op_tnl_4')
// (6, 5, 'neigh_op_lft_4')
// (6, 6, 'neigh_op_bnl_4')

wire n157;
// (4, 4, 'neigh_op_tnr_5')
// (4, 5, 'neigh_op_rgt_5')
// (4, 6, 'neigh_op_bnr_5')
// (5, 4, 'neigh_op_top_5')
// (5, 5, 'local_g0_5')
// (5, 5, 'local_g1_5')
// (5, 5, 'lutff_3/in_2')
// (5, 5, 'lutff_5/out')
// (5, 5, 'lutff_6/in_0')
// (5, 6, 'neigh_op_bot_5')
// (6, 4, 'neigh_op_tnl_5')
// (6, 5, 'neigh_op_lft_5')
// (6, 6, 'neigh_op_bnl_5')

wire n158;
// (4, 4, 'neigh_op_tnr_6')
// (4, 5, 'neigh_op_rgt_6')
// (4, 6, 'neigh_op_bnr_6')
// (5, 4, 'neigh_op_top_6')
// (5, 5, 'lutff_6/out')
// (5, 5, 'sp4_r_v_b_45')
// (5, 6, 'neigh_op_bot_6')
// (5, 6, 'sp4_r_v_b_32')
// (5, 7, 'sp4_r_v_b_21')
// (5, 8, 'sp4_r_v_b_8')
// (6, 4, 'local_g3_6')
// (6, 4, 'lutff_2/in_1')
// (6, 4, 'neigh_op_tnl_6')
// (6, 4, 'sp4_h_r_1')
// (6, 4, 'sp4_v_t_45')
// (6, 5, 'neigh_op_lft_6')
// (6, 5, 'sp4_v_b_45')
// (6, 6, 'neigh_op_bnl_6')
// (6, 6, 'sp4_v_b_32')
// (6, 7, 'sp4_v_b_21')
// (6, 8, 'sp4_v_b_8')
// (7, 4, 'local_g0_4')
// (7, 4, 'local_g1_4')
// (7, 4, 'lutff_3/in_3')
// (7, 4, 'lutff_4/in_3')
// (7, 4, 'sp4_h_r_12')
// (8, 4, 'sp4_h_r_25')
// (9, 4, 'sp4_h_r_36')
// (10, 4, 'sp4_h_l_36')

reg n159 = 0;
// (4, 4, 'neigh_op_tnr_7')
// (4, 5, 'neigh_op_rgt_7')
// (4, 6, 'neigh_op_bnr_7')
// (5, 4, 'neigh_op_top_7')
// (5, 5, 'local_g0_7')
// (5, 5, 'lutff_2/in_3')
// (5, 5, 'lutff_7/out')
// (5, 6, 'neigh_op_bot_7')
// (6, 4, 'neigh_op_tnl_7')
// (6, 5, 'neigh_op_lft_7')
// (6, 6, 'neigh_op_bnl_7')

wire n160;
// (4, 4, 'sp4_h_r_4')
// (5, 3, 'neigh_op_tnr_6')
// (5, 4, 'neigh_op_rgt_6')
// (5, 4, 'sp4_h_r_17')
// (5, 5, 'neigh_op_bnr_6')
// (6, 3, 'neigh_op_top_6')
// (6, 4, 'local_g0_6')
// (6, 4, 'lutff_4/in_2')
// (6, 4, 'lutff_6/out')
// (6, 4, 'sp4_h_r_28')
// (6, 5, 'neigh_op_bot_6')
// (7, 3, 'local_g2_6')
// (7, 3, 'lutff_3/in_1')
// (7, 3, 'lutff_4/in_2')
// (7, 3, 'neigh_op_tnl_6')
// (7, 4, 'local_g2_1')
// (7, 4, 'lutff_0/in_3')
// (7, 4, 'neigh_op_lft_6')
// (7, 4, 'sp4_h_r_41')
// (7, 5, 'neigh_op_bnl_6')
// (8, 4, 'sp4_h_l_41')

wire n161;
// (4, 4, 'sp4_h_r_8')
// (5, 3, 'neigh_op_tnr_0')
// (5, 4, 'neigh_op_rgt_0')
// (5, 4, 'sp4_h_r_21')
// (5, 4, 'sp4_h_r_5')
// (5, 5, 'neigh_op_bnr_0')
// (6, 3, 'neigh_op_top_0')
// (6, 4, 'lutff_0/out')
// (6, 4, 'sp4_h_r_16')
// (6, 4, 'sp4_h_r_32')
// (6, 5, 'neigh_op_bot_0')
// (7, 1, 'sp4_r_v_b_45')
// (7, 2, 'sp4_r_v_b_32')
// (7, 3, 'local_g2_0')
// (7, 3, 'local_g3_0')
// (7, 3, 'lutff_3/in_3')
// (7, 3, 'lutff_4/in_1')
// (7, 3, 'neigh_op_tnl_0')
// (7, 3, 'sp4_r_v_b_21')
// (7, 4, 'neigh_op_lft_0')
// (7, 4, 'sp4_h_r_29')
// (7, 4, 'sp4_h_r_45')
// (7, 4, 'sp4_r_v_b_8')
// (7, 5, 'neigh_op_bnl_0')
// (8, 0, 'span4_vert_45')
// (8, 1, 'sp4_r_v_b_46')
// (8, 1, 'sp4_v_b_45')
// (8, 2, 'sp4_r_v_b_35')
// (8, 2, 'sp4_v_b_32')
// (8, 3, 'local_g1_5')
// (8, 3, 'local_g3_6')
// (8, 3, 'lutff_0/in_3')
// (8, 3, 'lutff_5/in_1')
// (8, 3, 'sp4_r_v_b_22')
// (8, 3, 'sp4_v_b_21')
// (8, 4, 'sp4_h_l_45')
// (8, 4, 'sp4_h_r_40')
// (8, 4, 'sp4_r_v_b_11')
// (8, 4, 'sp4_v_b_8')
// (9, 0, 'span4_vert_46')
// (9, 1, 'sp4_v_b_46')
// (9, 2, 'sp4_v_b_35')
// (9, 3, 'sp4_v_b_22')
// (9, 4, 'sp4_h_l_40')
// (9, 4, 'sp4_v_b_11')

reg n162 = 0;
// (4, 4, 'sp4_r_v_b_45')
// (4, 5, 'sp4_r_v_b_32')
// (4, 6, 'neigh_op_tnr_4')
// (4, 6, 'sp4_r_v_b_21')
// (4, 7, 'neigh_op_rgt_4')
// (4, 7, 'sp4_r_v_b_8')
// (4, 8, 'neigh_op_bnr_4')
// (5, 3, 'sp4_v_t_45')
// (5, 4, 'sp4_v_b_45')
// (5, 5, 'sp4_v_b_32')
// (5, 6, 'local_g0_5')
// (5, 6, 'lutff_5/in_0')
// (5, 6, 'neigh_op_top_4')
// (5, 6, 'sp4_v_b_21')
// (5, 7, 'lutff_4/out')
// (5, 7, 'sp4_v_b_8')
// (5, 8, 'neigh_op_bot_4')
// (6, 6, 'neigh_op_tnl_4')
// (6, 7, 'neigh_op_lft_4')
// (6, 8, 'neigh_op_bnl_4')

wire n163;
// (4, 5, 'neigh_op_tnr_0')
// (4, 5, 'sp4_r_v_b_45')
// (4, 6, 'neigh_op_rgt_0')
// (4, 6, 'sp4_r_v_b_32')
// (4, 7, 'neigh_op_bnr_0')
// (4, 7, 'sp4_r_v_b_21')
// (4, 8, 'sp4_r_v_b_8')
// (5, 4, 'sp4_v_t_45')
// (5, 5, 'neigh_op_top_0')
// (5, 5, 'sp4_v_b_45')
// (5, 6, 'local_g1_0')
// (5, 6, 'lutff_0/out')
// (5, 6, 'lutff_3/in_2')
// (5, 6, 'sp4_v_b_32')
// (5, 7, 'local_g0_0')
// (5, 7, 'lutff_4/in_0')
// (5, 7, 'neigh_op_bot_0')
// (5, 7, 'sp4_v_b_21')
// (5, 8, 'local_g0_0')
// (5, 8, 'lutff_6/in_2')
// (5, 8, 'sp4_v_b_8')
// (6, 5, 'neigh_op_tnl_0')
// (6, 6, 'neigh_op_lft_0')
// (6, 7, 'neigh_op_bnl_0')

reg n164 = 0;
// (4, 5, 'neigh_op_tnr_3')
// (4, 6, 'neigh_op_rgt_3')
// (4, 7, 'neigh_op_bnr_3')
// (5, 5, 'neigh_op_top_3')
// (5, 6, 'local_g1_3')
// (5, 6, 'lutff_2/in_2')
// (5, 6, 'lutff_3/out')
// (5, 7, 'neigh_op_bot_3')
// (6, 5, 'neigh_op_tnl_3')
// (6, 6, 'neigh_op_lft_3')
// (6, 7, 'neigh_op_bnl_3')

reg n165 = 0;
// (4, 5, 'neigh_op_tnr_4')
// (4, 6, 'neigh_op_rgt_4')
// (4, 7, 'neigh_op_bnr_4')
// (5, 5, 'local_g1_4')
// (5, 5, 'lutff_4/in_3')
// (5, 5, 'neigh_op_top_4')
// (5, 6, 'local_g1_4')
// (5, 6, 'lutff_4/out')
// (5, 6, 'lutff_7/in_0')
// (5, 7, 'neigh_op_bot_4')
// (6, 5, 'neigh_op_tnl_4')
// (6, 6, 'neigh_op_lft_4')
// (6, 7, 'neigh_op_bnl_4')

reg n166 = 0;
// (4, 5, 'neigh_op_tnr_5')
// (4, 6, 'neigh_op_rgt_5')
// (4, 7, 'neigh_op_bnr_5')
// (5, 5, 'neigh_op_top_5')
// (5, 6, 'local_g1_5')
// (5, 6, 'lutff_4/in_0')
// (5, 6, 'lutff_5/out')
// (5, 7, 'neigh_op_bot_5')
// (6, 5, 'neigh_op_tnl_5')
// (6, 6, 'neigh_op_lft_5')
// (6, 7, 'neigh_op_bnl_5')

reg n167 = 0;
// (4, 5, 'neigh_op_tnr_6')
// (4, 6, 'neigh_op_rgt_6')
// (4, 7, 'neigh_op_bnr_6')
// (5, 0, 'span12_vert_23')
// (5, 1, 'sp12_v_b_23')
// (5, 2, 'sp12_v_b_20')
// (5, 3, 'sp12_v_b_19')
// (5, 4, 'sp12_v_b_16')
// (5, 4, 'sp4_r_v_b_37')
// (5, 5, 'neigh_op_top_6')
// (5, 5, 'sp12_v_b_15')
// (5, 5, 'sp4_r_v_b_24')
// (5, 6, 'lutff_6/out')
// (5, 6, 'sp12_v_b_12')
// (5, 6, 'sp4_r_v_b_13')
// (5, 7, 'neigh_op_bot_6')
// (5, 7, 'sp12_v_b_11')
// (5, 7, 'sp4_r_v_b_0')
// (5, 8, 'sp12_v_b_8')
// (5, 8, 'sp4_r_v_b_37')
// (5, 9, 'sp12_v_b_7')
// (5, 9, 'sp4_r_v_b_24')
// (5, 10, 'sp12_v_b_4')
// (5, 10, 'sp4_r_v_b_13')
// (5, 11, 'sp12_v_b_3')
// (5, 11, 'sp4_r_v_b_0')
// (5, 12, 'local_g2_0')
// (5, 12, 'lutff_0/in_0')
// (5, 12, 'sp12_h_r_0')
// (5, 12, 'sp12_v_b_0')
// (6, 3, 'sp4_v_t_37')
// (6, 4, 'sp4_v_b_37')
// (6, 5, 'neigh_op_tnl_6')
// (6, 5, 'sp4_v_b_24')
// (6, 6, 'local_g0_6')
// (6, 6, 'lutff_2/in_0')
// (6, 6, 'neigh_op_lft_6')
// (6, 6, 'sp4_v_b_13')
// (6, 7, 'neigh_op_bnl_6')
// (6, 7, 'sp4_v_b_0')
// (6, 7, 'sp4_v_t_37')
// (6, 8, 'sp4_v_b_37')
// (6, 9, 'sp4_v_b_24')
// (6, 10, 'sp4_v_b_13')
// (6, 11, 'sp4_h_r_6')
// (6, 11, 'sp4_v_b_0')
// (6, 12, 'sp12_h_r_3')
// (7, 11, 'local_g0_3')
// (7, 11, 'lutff_1/in_2')
// (7, 11, 'sp4_h_r_19')
// (7, 12, 'local_g1_4')
// (7, 12, 'lutff_5/in_2')
// (7, 12, 'sp12_h_r_4')
// (8, 11, 'sp4_h_r_30')
// (8, 12, 'sp12_h_r_7')
// (9, 11, 'sp4_h_r_43')
// (9, 12, 'sp12_h_r_8')
// (10, 11, 'sp4_h_l_43')
// (10, 12, 'sp12_h_r_11')
// (11, 12, 'sp12_h_r_12')
// (12, 12, 'sp12_h_r_15')
// (13, 12, 'span12_horz_15')

reg n168 = 0;
// (4, 5, 'neigh_op_tnr_7')
// (4, 5, 'sp4_r_v_b_43')
// (4, 6, 'neigh_op_rgt_7')
// (4, 6, 'sp4_r_v_b_30')
// (4, 7, 'neigh_op_bnr_7')
// (4, 7, 'sp4_r_v_b_19')
// (4, 8, 'sp4_r_v_b_6')
// (4, 9, 'sp4_r_v_b_44')
// (4, 10, 'sp4_r_v_b_33')
// (4, 11, 'sp4_r_v_b_20')
// (4, 12, 'sp4_r_v_b_9')
// (5, 4, 'sp4_v_t_43')
// (5, 5, 'neigh_op_top_7')
// (5, 5, 'sp4_r_v_b_42')
// (5, 5, 'sp4_v_b_43')
// (5, 6, 'lutff_7/out')
// (5, 6, 'sp4_r_v_b_31')
// (5, 6, 'sp4_v_b_30')
// (5, 7, 'neigh_op_bot_7')
// (5, 7, 'sp4_r_v_b_18')
// (5, 7, 'sp4_v_b_19')
// (5, 8, 'sp4_r_v_b_7')
// (5, 8, 'sp4_v_b_6')
// (5, 8, 'sp4_v_t_44')
// (5, 9, 'sp4_r_v_b_38')
// (5, 9, 'sp4_v_b_44')
// (5, 10, 'sp4_r_v_b_27')
// (5, 10, 'sp4_v_b_33')
// (5, 11, 'sp4_r_v_b_14')
// (5, 11, 'sp4_v_b_20')
// (5, 12, 'local_g0_1')
// (5, 12, 'lutff_1/in_0')
// (5, 12, 'sp4_r_v_b_3')
// (5, 12, 'sp4_v_b_9')
// (6, 4, 'sp4_v_t_42')
// (6, 5, 'neigh_op_tnl_7')
// (6, 5, 'sp4_v_b_42')
// (6, 6, 'local_g0_7')
// (6, 6, 'lutff_5/in_0')
// (6, 6, 'neigh_op_lft_7')
// (6, 6, 'sp4_v_b_31')
// (6, 7, 'neigh_op_bnl_7')
// (6, 7, 'sp4_v_b_18')
// (6, 8, 'sp4_v_b_7')
// (6, 8, 'sp4_v_t_38')
// (6, 9, 'sp4_v_b_38')
// (6, 10, 'sp4_v_b_27')
// (6, 11, 'local_g1_6')
// (6, 11, 'lutff_1/in_2')
// (6, 11, 'sp4_v_b_14')
// (6, 12, 'local_g0_1')
// (6, 12, 'lutff_5/in_2')
// (6, 12, 'sp4_h_r_9')
// (6, 12, 'sp4_v_b_3')
// (7, 12, 'sp4_h_r_20')
// (8, 12, 'sp4_h_r_33')
// (9, 12, 'sp4_h_r_44')
// (10, 12, 'sp4_h_l_44')

wire n169;
// (4, 5, 'sp12_h_r_1')
// (5, 5, 'sp12_h_r_2')
// (6, 4, 'neigh_op_tnr_7')
// (6, 5, 'neigh_op_rgt_7')
// (6, 5, 'sp12_h_r_5')
// (6, 6, 'neigh_op_bnr_7')
// (7, 4, 'neigh_op_top_7')
// (7, 5, 'lutff_7/out')
// (7, 5, 'sp12_h_r_6')
// (7, 6, 'neigh_op_bot_7')
// (8, 4, 'neigh_op_tnl_7')
// (8, 5, 'local_g1_1')
// (8, 5, 'lutff_5/in_3')
// (8, 5, 'neigh_op_lft_7')
// (8, 5, 'sp12_h_r_9')
// (8, 6, 'neigh_op_bnl_7')
// (9, 5, 'sp12_h_r_10')
// (10, 5, 'sp12_h_r_13')
// (11, 5, 'sp12_h_r_14')
// (12, 5, 'sp12_h_r_17')
// (13, 5, 'span12_horz_17')

wire n170;
// (4, 5, 'sp4_h_r_5')
// (5, 5, 'sp4_h_r_16')
// (6, 4, 'neigh_op_tnr_4')
// (6, 5, 'neigh_op_rgt_4')
// (6, 5, 'sp4_h_r_29')
// (6, 6, 'neigh_op_bnr_4')
// (7, 4, 'neigh_op_top_4')
// (7, 5, 'local_g2_0')
// (7, 5, 'lutff_4/out')
// (7, 5, 'lutff_5/in_3')
// (7, 5, 'sp4_h_r_40')
// (7, 6, 'neigh_op_bot_4')
// (8, 4, 'neigh_op_tnl_4')
// (8, 5, 'local_g1_4')
// (8, 5, 'lutff_3/in_2')
// (8, 5, 'neigh_op_lft_4')
// (8, 5, 'sp4_h_l_40')
// (8, 6, 'neigh_op_bnl_4')

wire n171;
// (4, 5, 'sp4_h_r_9')
// (5, 5, 'sp4_h_r_20')
// (6, 5, 'sp4_h_r_33')
// (7, 2, 'neigh_op_tnr_6')
// (7, 2, 'sp4_r_v_b_41')
// (7, 3, 'neigh_op_rgt_6')
// (7, 3, 'sp4_r_v_b_28')
// (7, 4, 'neigh_op_bnr_6')
// (7, 4, 'sp4_r_v_b_17')
// (7, 5, 'local_g2_4')
// (7, 5, 'lutff_3/in_1')
// (7, 5, 'sp4_h_r_44')
// (7, 5, 'sp4_r_v_b_4')
// (8, 1, 'sp4_v_t_41')
// (8, 2, 'neigh_op_top_6')
// (8, 2, 'sp4_v_b_41')
// (8, 3, 'lutff_6/out')
// (8, 3, 'sp4_v_b_28')
// (8, 4, 'local_g0_6')
// (8, 4, 'lutff_3/in_1')
// (8, 4, 'neigh_op_bot_6')
// (8, 4, 'sp4_v_b_17')
// (8, 5, 'local_g0_4')
// (8, 5, 'lutff_4/in_2')
// (8, 5, 'sp4_h_l_44')
// (8, 5, 'sp4_v_b_4')
// (9, 2, 'neigh_op_tnl_6')
// (9, 3, 'neigh_op_lft_6')
// (9, 4, 'neigh_op_bnl_6')

reg n172 = 0;
// (4, 5, 'sp4_r_v_b_37')
// (4, 6, 'sp4_r_v_b_24')
// (4, 7, 'neigh_op_tnr_0')
// (4, 7, 'sp4_r_v_b_13')
// (4, 8, 'neigh_op_rgt_0')
// (4, 8, 'sp4_r_v_b_0')
// (4, 9, 'neigh_op_bnr_0')
// (5, 4, 'sp4_v_t_37')
// (5, 5, 'sp4_v_b_37')
// (5, 6, 'local_g3_0')
// (5, 6, 'lutff_0/in_3')
// (5, 6, 'lutff_2/in_1')
// (5, 6, 'sp4_v_b_24')
// (5, 7, 'neigh_op_top_0')
// (5, 7, 'sp4_v_b_13')
// (5, 8, 'lutff_0/out')
// (5, 8, 'sp4_v_b_0')
// (5, 9, 'neigh_op_bot_0')
// (6, 7, 'neigh_op_tnl_0')
// (6, 8, 'neigh_op_lft_0')
// (6, 9, 'neigh_op_bnl_0')

wire n173;
// (4, 5, 'sp4_r_v_b_38')
// (4, 6, 'local_g0_3')
// (4, 6, 'lutff_2/in_1')
// (4, 6, 'sp4_r_v_b_27')
// (4, 7, 'sp4_r_v_b_14')
// (4, 8, 'sp4_r_v_b_3')
// (5, 4, 'sp4_h_r_3')
// (5, 4, 'sp4_v_t_38')
// (5, 5, 'sp4_v_b_38')
// (5, 6, 'sp4_v_b_27')
// (5, 7, 'sp4_v_b_14')
// (5, 8, 'sp4_v_b_3')
// (6, 4, 'sp4_h_r_14')
// (7, 3, 'neigh_op_tnr_3')
// (7, 4, 'neigh_op_rgt_3')
// (7, 4, 'sp4_h_r_27')
// (7, 5, 'neigh_op_bnr_3')
// (8, 3, 'neigh_op_top_3')
// (8, 4, 'lutff_3/out')
// (8, 4, 'sp4_h_r_38')
// (8, 5, 'neigh_op_bot_3')
// (9, 3, 'neigh_op_tnl_3')
// (9, 4, 'neigh_op_lft_3')
// (9, 4, 'sp4_h_l_38')
// (9, 5, 'neigh_op_bnl_3')

reg n174 = 0;
// (4, 6, 'neigh_op_tnr_5')
// (4, 7, 'neigh_op_rgt_5')
// (4, 8, 'neigh_op_bnr_5')
// (5, 6, 'neigh_op_top_5')
// (5, 7, 'lutff_5/out')
// (5, 8, 'local_g1_5')
// (5, 8, 'lutff_4/in_0')
// (5, 8, 'neigh_op_bot_5')
// (6, 6, 'neigh_op_tnl_5')
// (6, 7, 'neigh_op_lft_5')
// (6, 8, 'neigh_op_bnl_5')

wire n175;
// (4, 6, 'sp4_h_r_4')
// (5, 6, 'local_g0_1')
// (5, 6, 'lutff_0/in_1')
// (5, 6, 'sp4_h_r_17')
// (6, 6, 'sp4_h_r_28')
// (7, 3, 'neigh_op_tnr_6')
// (7, 3, 'sp4_r_v_b_41')
// (7, 4, 'neigh_op_rgt_6')
// (7, 4, 'sp4_r_v_b_28')
// (7, 5, 'local_g1_6')
// (7, 5, 'lutff_3/in_0')
// (7, 5, 'lutff_6/in_3')
// (7, 5, 'neigh_op_bnr_6')
// (7, 5, 'sp4_r_v_b_17')
// (7, 6, 'sp4_h_r_41')
// (7, 6, 'sp4_r_v_b_4')
// (8, 2, 'sp4_v_t_41')
// (8, 3, 'neigh_op_top_6')
// (8, 3, 'sp4_v_b_41')
// (8, 4, 'lutff_6/out')
// (8, 4, 'sp4_v_b_28')
// (8, 5, 'local_g0_6')
// (8, 5, 'lutff_4/in_0')
// (8, 5, 'neigh_op_bot_6')
// (8, 5, 'sp4_v_b_17')
// (8, 6, 'sp4_h_l_41')
// (8, 6, 'sp4_v_b_4')
// (9, 3, 'neigh_op_tnl_6')
// (9, 4, 'neigh_op_lft_6')
// (9, 5, 'neigh_op_bnl_6')

wire n176;
// (4, 6, 'sp4_h_r_7')
// (5, 6, 'local_g0_2')
// (5, 6, 'lutff_3/in_3')
// (5, 6, 'sp4_h_r_18')
// (6, 6, 'sp4_h_r_31')
// (7, 6, 'neigh_op_tnr_2')
// (7, 6, 'sp4_h_r_42')
// (7, 7, 'neigh_op_rgt_2')
// (7, 7, 'sp4_r_v_b_36')
// (7, 8, 'neigh_op_bnr_2')
// (7, 8, 'sp4_r_v_b_25')
// (7, 9, 'sp4_r_v_b_12')
// (7, 10, 'sp4_r_v_b_1')
// (7, 11, 'local_g3_4')
// (7, 11, 'lutff_4/in_3')
// (7, 11, 'sp4_r_v_b_44')
// (7, 12, 'sp4_r_v_b_33')
// (7, 13, 'sp4_r_v_b_20')
// (7, 14, 'sp4_r_v_b_9')
// (8, 5, 'sp4_r_v_b_45')
// (8, 6, 'neigh_op_top_2')
// (8, 6, 'sp4_h_l_42')
// (8, 6, 'sp4_r_v_b_32')
// (8, 6, 'sp4_v_t_36')
// (8, 7, 'lutff_2/out')
// (8, 7, 'sp4_r_v_b_21')
// (8, 7, 'sp4_v_b_36')
// (8, 8, 'neigh_op_bot_2')
// (8, 8, 'sp4_r_v_b_8')
// (8, 8, 'sp4_v_b_25')
// (8, 9, 'local_g1_4')
// (8, 9, 'lutff_0/in_3')
// (8, 9, 'lutff_2/in_3')
// (8, 9, 'lutff_6/in_3')
// (8, 9, 'sp4_r_v_b_46')
// (8, 9, 'sp4_v_b_12')
// (8, 10, 'local_g0_1')
// (8, 10, 'lutff_1/in_2')
// (8, 10, 'sp4_r_v_b_35')
// (8, 10, 'sp4_v_b_1')
// (8, 10, 'sp4_v_t_44')
// (8, 11, 'local_g3_4')
// (8, 11, 'lutff_2/in_3')
// (8, 11, 'sp4_r_v_b_22')
// (8, 11, 'sp4_v_b_44')
// (8, 12, 'local_g2_1')
// (8, 12, 'lutff_0/in_3')
// (8, 12, 'sp4_r_v_b_11')
// (8, 12, 'sp4_v_b_33')
// (8, 13, 'sp4_v_b_20')
// (8, 14, 'sp4_v_b_9')
// (9, 4, 'sp4_v_t_45')
// (9, 5, 'sp4_v_b_45')
// (9, 6, 'neigh_op_tnl_2')
// (9, 6, 'sp4_v_b_32')
// (9, 7, 'neigh_op_lft_2')
// (9, 7, 'sp4_v_b_21')
// (9, 8, 'neigh_op_bnl_2')
// (9, 8, 'sp4_v_b_8')
// (9, 8, 'sp4_v_t_46')
// (9, 9, 'sp4_v_b_46')
// (9, 10, 'sp4_v_b_35')
// (9, 11, 'sp4_v_b_22')
// (9, 12, 'local_g0_3')
// (9, 12, 'lutff_6/in_3')
// (9, 12, 'sp4_v_b_11')

reg n177 = 0;
// (4, 7, 'neigh_op_tnr_1')
// (4, 8, 'neigh_op_rgt_1')
// (4, 9, 'neigh_op_bnr_1')
// (5, 7, 'neigh_op_top_1')
// (5, 8, 'local_g1_1')
// (5, 8, 'lutff_0/in_0')
// (5, 8, 'lutff_1/out')
// (5, 9, 'neigh_op_bot_1')
// (6, 7, 'neigh_op_tnl_1')
// (6, 8, 'neigh_op_lft_1')
// (6, 9, 'neigh_op_bnl_1')

reg n178 = 0;
// (4, 7, 'neigh_op_tnr_2')
// (4, 8, 'neigh_op_rgt_2')
// (4, 9, 'neigh_op_bnr_2')
// (5, 7, 'neigh_op_top_2')
// (5, 8, 'local_g1_2')
// (5, 8, 'lutff_1/in_0')
// (5, 8, 'lutff_2/out')
// (5, 9, 'neigh_op_bot_2')
// (6, 7, 'neigh_op_tnl_2')
// (6, 8, 'neigh_op_lft_2')
// (6, 9, 'neigh_op_bnl_2')

reg n179 = 0;
// (4, 7, 'neigh_op_tnr_4')
// (4, 8, 'neigh_op_rgt_4')
// (4, 9, 'neigh_op_bnr_4')
// (5, 7, 'neigh_op_top_4')
// (5, 8, 'local_g1_4')
// (5, 8, 'lutff_4/out')
// (5, 8, 'lutff_5/in_0')
// (5, 9, 'neigh_op_bot_4')
// (6, 7, 'neigh_op_tnl_4')
// (6, 8, 'neigh_op_lft_4')
// (6, 9, 'neigh_op_bnl_4')

reg n180 = 0;
// (4, 7, 'neigh_op_tnr_5')
// (4, 8, 'neigh_op_rgt_5')
// (4, 9, 'neigh_op_bnr_5')
// (5, 1, 'sp12_v_t_22')
// (5, 2, 'sp12_v_b_22')
// (5, 3, 'sp12_v_b_21')
// (5, 4, 'sp12_v_b_18')
// (5, 5, 'local_g3_1')
// (5, 5, 'lutff_5/in_3')
// (5, 5, 'sp12_v_b_17')
// (5, 6, 'sp12_v_b_14')
// (5, 7, 'neigh_op_top_5')
// (5, 7, 'sp12_v_b_13')
// (5, 8, 'local_g2_5')
// (5, 8, 'lutff_3/in_0')
// (5, 8, 'lutff_5/out')
// (5, 8, 'sp12_v_b_10')
// (5, 9, 'neigh_op_bot_5')
// (5, 9, 'sp12_v_b_9')
// (5, 10, 'sp12_v_b_6')
// (5, 11, 'sp12_v_b_5')
// (5, 12, 'sp12_v_b_2')
// (5, 13, 'sp12_v_b_1')
// (6, 7, 'neigh_op_tnl_5')
// (6, 8, 'neigh_op_lft_5')
// (6, 9, 'neigh_op_bnl_5')

reg n181 = 0;
// (4, 7, 'neigh_op_tnr_6')
// (4, 8, 'neigh_op_rgt_6')
// (4, 9, 'neigh_op_bnr_6')
// (5, 7, 'neigh_op_top_6')
// (5, 8, 'local_g0_6')
// (5, 8, 'lutff_2/in_0')
// (5, 8, 'lutff_6/out')
// (5, 9, 'neigh_op_bot_6')
// (6, 7, 'neigh_op_tnl_6')
// (6, 8, 'neigh_op_lft_6')
// (6, 9, 'neigh_op_bnl_6')

reg n182 = 0;
// (4, 7, 'neigh_op_tnr_7')
// (4, 8, 'neigh_op_rgt_7')
// (4, 9, 'neigh_op_bnr_7')
// (5, 7, 'neigh_op_top_7')
// (5, 8, 'local_g0_7')
// (5, 8, 'lutff_6/in_3')
// (5, 8, 'lutff_7/out')
// (5, 9, 'neigh_op_bot_7')
// (6, 7, 'neigh_op_tnl_7')
// (6, 8, 'neigh_op_lft_7')
// (6, 9, 'neigh_op_bnl_7')

wire n183;
// (4, 7, 'sp4_h_r_10')
// (5, 6, 'neigh_op_tnr_1')
// (5, 7, 'neigh_op_rgt_1')
// (5, 7, 'sp4_h_r_23')
// (5, 8, 'neigh_op_bnr_1')
// (6, 6, 'neigh_op_top_1')
// (6, 7, 'local_g2_1')
// (6, 7, 'lutff_1/out')
// (6, 7, 'lutff_6/in_3')
// (6, 7, 'sp4_h_r_34')
// (6, 8, 'neigh_op_bot_1')
// (7, 4, 'sp4_r_v_b_41')
// (7, 5, 'sp4_r_v_b_28')
// (7, 6, 'neigh_op_tnl_1')
// (7, 6, 'sp4_r_v_b_17')
// (7, 7, 'local_g1_1')
// (7, 7, 'lutff_1/in_1')
// (7, 7, 'lutff_3/in_1')
// (7, 7, 'neigh_op_lft_1')
// (7, 7, 'sp4_h_r_47')
// (7, 7, 'sp4_r_v_b_4')
// (7, 8, 'neigh_op_bnl_1')
// (8, 3, 'sp4_v_t_41')
// (8, 4, 'sp4_v_b_41')
// (8, 5, 'sp4_v_b_28')
// (8, 6, 'local_g0_1')
// (8, 6, 'local_g1_1')
// (8, 6, 'lutff_0/in_2')
// (8, 6, 'lutff_3/in_2')
// (8, 6, 'sp4_v_b_17')
// (8, 7, 'sp4_h_l_47')
// (8, 7, 'sp4_v_b_4')

wire n184;
// (4, 7, 'sp4_h_r_6')
// (5, 6, 'neigh_op_tnr_7')
// (5, 7, 'neigh_op_rgt_7')
// (5, 7, 'sp4_h_r_19')
// (5, 8, 'neigh_op_bnr_7')
// (6, 6, 'neigh_op_top_7')
// (6, 7, 'local_g3_7')
// (6, 7, 'lutff_6/in_2')
// (6, 7, 'lutff_7/out')
// (6, 7, 'sp4_h_r_30')
// (6, 8, 'neigh_op_bot_7')
// (7, 4, 'sp4_r_v_b_43')
// (7, 5, 'sp4_r_v_b_30')
// (7, 6, 'neigh_op_tnl_7')
// (7, 6, 'sp4_r_v_b_19')
// (7, 7, 'local_g0_7')
// (7, 7, 'lutff_1/in_0')
// (7, 7, 'lutff_3/in_0')
// (7, 7, 'neigh_op_lft_7')
// (7, 7, 'sp4_h_r_43')
// (7, 7, 'sp4_r_v_b_6')
// (7, 8, 'neigh_op_bnl_7')
// (8, 3, 'sp4_v_t_43')
// (8, 4, 'sp4_v_b_43')
// (8, 5, 'sp4_v_b_30')
// (8, 6, 'local_g0_3')
// (8, 6, 'lutff_1/in_2')
// (8, 6, 'lutff_7/in_2')
// (8, 6, 'sp4_v_b_19')
// (8, 7, 'sp4_h_l_43')
// (8, 7, 'sp4_v_b_6')

reg n185 = 0;
// (4, 8, 'neigh_op_tnr_0')
// (4, 9, 'neigh_op_rgt_0')
// (4, 10, 'neigh_op_bnr_0')
// (5, 8, 'neigh_op_top_0')
// (5, 9, 'local_g0_0')
// (5, 9, 'lutff_0/out')
// (5, 9, 'lutff_6/in_0')
// (5, 10, 'neigh_op_bot_0')
// (6, 8, 'neigh_op_tnl_0')
// (6, 9, 'neigh_op_lft_0')
// (6, 10, 'neigh_op_bnl_0')

reg n186 = 0;
// (4, 8, 'neigh_op_tnr_1')
// (4, 9, 'neigh_op_rgt_1')
// (4, 10, 'neigh_op_bnr_1')
// (5, 8, 'neigh_op_top_1')
// (5, 9, 'local_g1_1')
// (5, 9, 'lutff_1/out')
// (5, 9, 'lutff_2/in_0')
// (5, 10, 'neigh_op_bot_1')
// (6, 8, 'neigh_op_tnl_1')
// (6, 9, 'neigh_op_lft_1')
// (6, 10, 'neigh_op_bnl_1')

reg n187 = 0;
// (4, 8, 'neigh_op_tnr_2')
// (4, 9, 'neigh_op_rgt_2')
// (4, 10, 'neigh_op_bnr_2')
// (5, 8, 'neigh_op_top_2')
// (5, 9, 'local_g0_2')
// (5, 9, 'lutff_2/out')
// (5, 9, 'lutff_7/in_1')
// (5, 9, 'sp4_h_r_4')
// (5, 10, 'neigh_op_bot_2')
// (6, 8, 'neigh_op_tnl_2')
// (6, 9, 'local_g0_1')
// (6, 9, 'lutff_2/in_1')
// (6, 9, 'neigh_op_lft_2')
// (6, 9, 'sp4_h_r_17')
// (6, 10, 'neigh_op_bnl_2')
// (7, 9, 'sp4_h_r_28')
// (8, 9, 'sp4_h_r_41')
// (9, 9, 'sp4_h_l_41')

reg n188 = 0;
// (4, 8, 'neigh_op_tnr_3')
// (4, 9, 'local_g3_3')
// (4, 9, 'lutff_3/in_1')
// (4, 9, 'neigh_op_rgt_3')
// (4, 10, 'neigh_op_bnr_3')
// (5, 8, 'neigh_op_top_3')
// (5, 9, 'lutff_3/out')
// (5, 10, 'neigh_op_bot_3')
// (6, 8, 'neigh_op_tnl_3')
// (6, 9, 'local_g1_3')
// (6, 9, 'lutff_2/in_0')
// (6, 9, 'neigh_op_lft_3')
// (6, 10, 'neigh_op_bnl_3')

reg n189 = 0;
// (4, 8, 'neigh_op_tnr_4')
// (4, 9, 'neigh_op_rgt_4')
// (4, 10, 'neigh_op_bnr_4')
// (5, 8, 'neigh_op_top_4')
// (5, 9, 'lutff_4/out')
// (5, 9, 'sp4_h_r_8')
// (5, 10, 'neigh_op_bot_4')
// (6, 8, 'neigh_op_tnl_4')
// (6, 9, 'neigh_op_lft_4')
// (6, 9, 'sp4_h_r_21')
// (6, 10, 'neigh_op_bnl_4')
// (7, 9, 'local_g2_0')
// (7, 9, 'lutff_4/in_0')
// (7, 9, 'sp4_h_r_32')
// (8, 9, 'sp4_h_r_45')
// (9, 9, 'sp4_h_l_45')

reg n190 = 0;
// (4, 8, 'neigh_op_tnr_6')
// (4, 9, 'neigh_op_rgt_6')
// (4, 10, 'neigh_op_bnr_6')
// (5, 8, 'neigh_op_top_6')
// (5, 8, 'sp4_r_v_b_40')
// (5, 9, 'local_g0_5')
// (5, 9, 'lutff_3/in_0')
// (5, 9, 'lutff_6/out')
// (5, 9, 'sp4_r_v_b_29')
// (5, 10, 'neigh_op_bot_6')
// (5, 10, 'sp4_r_v_b_16')
// (5, 11, 'sp4_r_v_b_5')
// (6, 7, 'sp4_v_t_40')
// (6, 8, 'neigh_op_tnl_6')
// (6, 8, 'sp4_v_b_40')
// (6, 9, 'neigh_op_lft_6')
// (6, 9, 'sp4_v_b_29')
// (6, 10, 'neigh_op_bnl_6')
// (6, 10, 'sp4_v_b_16')
// (6, 11, 'sp4_v_b_5')

reg n191 = 0;
// (4, 8, 'neigh_op_tnr_7')
// (4, 9, 'neigh_op_rgt_7')
// (4, 10, 'neigh_op_bnr_7')
// (5, 8, 'neigh_op_top_7')
// (5, 9, 'local_g1_7')
// (5, 9, 'lutff_0/in_0')
// (5, 9, 'lutff_7/out')
// (5, 10, 'neigh_op_bot_7')
// (6, 8, 'neigh_op_tnl_7')
// (6, 9, 'neigh_op_lft_7')
// (6, 10, 'neigh_op_bnl_7')

wire n192;
// (4, 8, 'sp4_h_r_6')
// (5, 7, 'neigh_op_tnr_7')
// (5, 8, 'neigh_op_rgt_7')
// (5, 8, 'sp4_h_r_19')
// (5, 9, 'neigh_op_bnr_7')
// (6, 7, 'local_g0_7')
// (6, 7, 'lutff_3/in_0')
// (6, 7, 'neigh_op_top_7')
// (6, 8, 'local_g0_7')
// (6, 8, 'lutff_4/in_3')
// (6, 8, 'lutff_7/out')
// (6, 8, 'sp4_h_r_30')
// (6, 9, 'neigh_op_bot_7')
// (7, 7, 'local_g2_7')
// (7, 7, 'lutff_4/in_1')
// (7, 7, 'neigh_op_tnl_7')
// (7, 8, 'local_g2_3')
// (7, 8, 'local_g3_3')
// (7, 8, 'lutff_2/in_3')
// (7, 8, 'lutff_4/in_0')
// (7, 8, 'neigh_op_lft_7')
// (7, 8, 'sp4_h_r_43')
// (7, 9, 'neigh_op_bnl_7')
// (8, 8, 'sp4_h_l_43')

wire n193;
// (4, 8, 'sp4_h_r_7')
// (5, 8, 'sp4_h_r_18')
// (6, 6, 'neigh_op_tnr_7')
// (6, 7, 'neigh_op_rgt_7')
// (6, 8, 'neigh_op_bnr_7')
// (6, 8, 'sp4_h_r_31')
// (7, 5, 'sp4_r_v_b_39')
// (7, 6, 'neigh_op_top_7')
// (7, 6, 'sp4_r_v_b_26')
// (7, 7, 'lutff_7/out')
// (7, 7, 'sp4_r_v_b_15')
// (7, 8, 'local_g1_2')
// (7, 8, 'local_g2_2')
// (7, 8, 'lutff_0/in_1')
// (7, 8, 'lutff_6/in_0')
// (7, 8, 'lutff_7/in_3')
// (7, 8, 'neigh_op_bot_7')
// (7, 8, 'sp4_h_r_42')
// (7, 8, 'sp4_r_v_b_2')
// (8, 4, 'sp4_v_t_39')
// (8, 5, 'sp4_v_b_39')
// (8, 6, 'local_g2_7')
// (8, 6, 'local_g3_7')
// (8, 6, 'lutff_2/in_1')
// (8, 6, 'lutff_4/in_3')
// (8, 6, 'lutff_5/in_1')
// (8, 6, 'lutff_6/in_3')
// (8, 6, 'neigh_op_tnl_7')
// (8, 6, 'sp4_v_b_26')
// (8, 7, 'local_g1_7')
// (8, 7, 'lutff_1/in_3')
// (8, 7, 'neigh_op_lft_7')
// (8, 7, 'sp4_v_b_15')
// (8, 8, 'neigh_op_bnl_7')
// (8, 8, 'sp4_h_l_42')
// (8, 8, 'sp4_v_b_2')

reg n194 = 0;
// (4, 8, 'sp4_r_v_b_45')
// (4, 9, 'sp4_r_v_b_32')
// (4, 10, 'neigh_op_tnr_4')
// (4, 10, 'sp4_r_v_b_21')
// (4, 11, 'neigh_op_rgt_4')
// (4, 11, 'sp4_r_v_b_8')
// (4, 12, 'neigh_op_bnr_4')
// (5, 7, 'sp4_v_t_45')
// (5, 8, 'sp4_v_b_45')
// (5, 9, 'sp4_v_b_32')
// (5, 10, 'local_g0_5')
// (5, 10, 'lutff_1/in_0')
// (5, 10, 'lutff_7/in_0')
// (5, 10, 'neigh_op_top_4')
// (5, 10, 'sp4_v_b_21')
// (5, 11, 'local_g1_4')
// (5, 11, 'lutff_4/out')
// (5, 11, 'lutff_5/in_0')
// (5, 11, 'lutff_7/in_0')
// (5, 11, 'sp4_v_b_8')
// (5, 12, 'neigh_op_bot_4')
// (6, 10, 'neigh_op_tnl_4')
// (6, 11, 'neigh_op_lft_4')
// (6, 12, 'neigh_op_bnl_4')

wire n195;
// (4, 9, 'neigh_op_tnr_1')
// (4, 10, 'neigh_op_rgt_1')
// (4, 11, 'neigh_op_bnr_1')
// (5, 9, 'neigh_op_top_1')
// (5, 10, 'local_g2_1')
// (5, 10, 'lutff_1/out')
// (5, 10, 'lutff_2/in_3')
// (5, 11, 'neigh_op_bot_1')
// (6, 9, 'neigh_op_tnl_1')
// (6, 10, 'neigh_op_lft_1')
// (6, 11, 'neigh_op_bnl_1')

wire n196;
// (4, 9, 'neigh_op_tnr_2')
// (4, 10, 'neigh_op_rgt_2')
// (4, 11, 'neigh_op_bnr_2')
// (5, 7, 'sp4_r_v_b_40')
// (5, 8, 'sp4_r_v_b_29')
// (5, 9, 'neigh_op_top_2')
// (5, 9, 'sp4_r_v_b_16')
// (5, 10, 'lutff_2/out')
// (5, 10, 'sp4_r_v_b_5')
// (5, 11, 'neigh_op_bot_2')
// (6, 6, 'sp4_v_t_40')
// (6, 7, 'sp4_v_b_40')
// (6, 8, 'local_g2_5')
// (6, 8, 'local_g3_5')
// (6, 8, 'lutff_2/in_0')
// (6, 8, 'lutff_3/in_0')
// (6, 8, 'lutff_5/in_0')
// (6, 8, 'lutff_7/in_1')
// (6, 8, 'sp4_v_b_29')
// (6, 9, 'local_g2_2')
// (6, 9, 'lutff_5/in_1')
// (6, 9, 'neigh_op_tnl_2')
// (6, 9, 'sp4_v_b_16')
// (6, 10, 'neigh_op_lft_2')
// (6, 10, 'sp4_v_b_5')
// (6, 11, 'neigh_op_bnl_2')

reg n197 = 0;
// (4, 9, 'neigh_op_tnr_4')
// (4, 10, 'neigh_op_rgt_4')
// (4, 11, 'neigh_op_bnr_4')
// (5, 9, 'neigh_op_top_4')
// (5, 10, 'local_g3_4')
// (5, 10, 'lutff_3/in_0')
// (5, 10, 'lutff_4/out')
// (5, 11, 'neigh_op_bot_4')
// (6, 9, 'neigh_op_tnl_4')
// (6, 10, 'neigh_op_lft_4')
// (6, 11, 'neigh_op_bnl_4')

reg n198 = 0;
// (4, 9, 'neigh_op_tnr_6')
// (4, 10, 'neigh_op_rgt_6')
// (4, 11, 'neigh_op_bnr_6')
// (5, 9, 'neigh_op_top_6')
// (5, 10, 'lutff_6/out')
// (5, 11, 'local_g0_6')
// (5, 11, 'lutff_2/in_0')
// (5, 11, 'neigh_op_bot_6')
// (6, 9, 'neigh_op_tnl_6')
// (6, 10, 'neigh_op_lft_6')
// (6, 11, 'neigh_op_bnl_6')

reg n199 = 0;
// (4, 9, 'neigh_op_tnr_7')
// (4, 10, 'neigh_op_rgt_7')
// (4, 11, 'neigh_op_bnr_7')
// (5, 9, 'neigh_op_top_7')
// (5, 10, 'local_g1_7')
// (5, 10, 'lutff_6/in_0')
// (5, 10, 'lutff_7/out')
// (5, 11, 'neigh_op_bot_7')
// (6, 9, 'neigh_op_tnl_7')
// (6, 10, 'neigh_op_lft_7')
// (6, 11, 'neigh_op_bnl_7')

wire n200;
// (4, 10, 'neigh_op_tnr_0')
// (4, 11, 'neigh_op_rgt_0')
// (4, 12, 'neigh_op_bnr_0')
// (5, 9, 'sp4_r_v_b_41')
// (5, 10, 'local_g0_4')
// (5, 10, 'lutff_1/in_3')
// (5, 10, 'neigh_op_top_0')
// (5, 10, 'sp4_r_v_b_28')
// (5, 11, 'lutff_0/out')
// (5, 11, 'sp4_r_v_b_17')
// (5, 12, 'neigh_op_bot_0')
// (5, 12, 'sp4_r_v_b_4')
// (6, 8, 'sp4_v_t_41')
// (6, 9, 'sp4_v_b_41')
// (6, 10, 'neigh_op_tnl_0')
// (6, 10, 'sp4_v_b_28')
// (6, 11, 'neigh_op_lft_0')
// (6, 11, 'sp4_v_b_17')
// (6, 12, 'neigh_op_bnl_0')
// (6, 12, 'sp4_v_b_4')

reg n201 = 0;
// (4, 10, 'neigh_op_tnr_1')
// (4, 11, 'neigh_op_rgt_1')
// (4, 12, 'neigh_op_bnr_1')
// (5, 10, 'neigh_op_top_1')
// (5, 11, 'local_g0_1')
// (5, 11, 'local_g1_1')
// (5, 11, 'lutff_0/in_1')
// (5, 11, 'lutff_1/out')
// (5, 11, 'lutff_5/in_1')
// (5, 12, 'neigh_op_bot_1')
// (6, 10, 'neigh_op_tnl_1')
// (6, 11, 'neigh_op_lft_1')
// (6, 12, 'neigh_op_bnl_1')

reg n202 = 0;
// (4, 10, 'neigh_op_tnr_2')
// (4, 11, 'neigh_op_rgt_2')
// (4, 12, 'neigh_op_bnr_2')
// (5, 10, 'neigh_op_top_2')
// (5, 11, 'local_g1_2')
// (5, 11, 'lutff_1/in_0')
// (5, 11, 'lutff_2/out')
// (5, 12, 'neigh_op_bot_2')
// (6, 10, 'neigh_op_tnl_2')
// (6, 11, 'neigh_op_lft_2')
// (6, 12, 'neigh_op_bnl_2')

reg n203 = 0;
// (4, 10, 'neigh_op_tnr_3')
// (4, 11, 'neigh_op_rgt_3')
// (4, 12, 'neigh_op_bnr_3')
// (5, 10, 'neigh_op_top_3')
// (5, 11, 'local_g1_3')
// (5, 11, 'lutff_3/out')
// (5, 11, 'lutff_4/in_0')
// (5, 12, 'neigh_op_bot_3')
// (6, 10, 'neigh_op_tnl_3')
// (6, 11, 'neigh_op_lft_3')
// (6, 12, 'neigh_op_bnl_3')

reg n204 = 0;
// (4, 10, 'neigh_op_tnr_5')
// (4, 11, 'local_g3_5')
// (4, 11, 'lutff_2/in_0')
// (4, 11, 'neigh_op_rgt_5')
// (4, 12, 'neigh_op_bnr_5')
// (5, 10, 'neigh_op_top_5')
// (5, 11, 'lutff_5/out')
// (5, 12, 'neigh_op_bot_5')
// (6, 10, 'neigh_op_tnl_5')
// (6, 11, 'neigh_op_lft_5')
// (6, 12, 'neigh_op_bnl_5')

reg n205 = 0;
// (4, 10, 'neigh_op_tnr_6')
// (4, 11, 'neigh_op_rgt_6')
// (4, 12, 'neigh_op_bnr_6')
// (5, 10, 'neigh_op_top_6')
// (5, 11, 'local_g1_6')
// (5, 11, 'lutff_3/in_0')
// (5, 11, 'lutff_6/out')
// (5, 12, 'neigh_op_bot_6')
// (6, 10, 'neigh_op_tnl_6')
// (6, 11, 'neigh_op_lft_6')
// (6, 12, 'neigh_op_bnl_6')

reg n206 = 0;
// (4, 10, 'neigh_op_tnr_7')
// (4, 11, 'neigh_op_rgt_7')
// (4, 12, 'neigh_op_bnr_7')
// (5, 10, 'neigh_op_top_7')
// (5, 11, 'local_g1_7')
// (5, 11, 'lutff_6/in_0')
// (5, 11, 'lutff_7/out')
// (5, 12, 'neigh_op_bot_7')
// (6, 10, 'neigh_op_tnl_7')
// (6, 11, 'neigh_op_lft_7')
// (6, 12, 'neigh_op_bnl_7')

reg n207 = 0;
// (4, 11, 'neigh_op_tnr_0')
// (4, 12, 'neigh_op_rgt_0')
// (4, 13, 'neigh_op_bnr_0')
// (5, 11, 'neigh_op_top_0')
// (5, 12, 'local_g0_0')
// (5, 12, 'lutff_0/out')
// (5, 12, 'lutff_4/in_0')
// (5, 13, 'neigh_op_bot_0')
// (6, 11, 'neigh_op_tnl_0')
// (6, 12, 'neigh_op_lft_0')
// (6, 13, 'neigh_op_bnl_0')

reg n208 = 0;
// (4, 11, 'neigh_op_tnr_1')
// (4, 12, 'local_g3_1')
// (4, 12, 'lutff_2/in_0')
// (4, 12, 'neigh_op_rgt_1')
// (4, 13, 'neigh_op_bnr_1')
// (5, 11, 'neigh_op_top_1')
// (5, 12, 'lutff_1/out')
// (5, 13, 'neigh_op_bot_1')
// (6, 11, 'neigh_op_tnl_1')
// (6, 12, 'neigh_op_lft_1')
// (6, 13, 'neigh_op_bnl_1')

reg n209 = 0;
// (4, 11, 'neigh_op_tnr_2')
// (4, 12, 'neigh_op_rgt_2')
// (4, 13, 'neigh_op_bnr_2')
// (5, 11, 'neigh_op_top_2')
// (5, 12, 'local_g3_2')
// (5, 12, 'lutff_2/out')
// (5, 12, 'lutff_3/in_0')
// (5, 13, 'neigh_op_bot_2')
// (6, 11, 'neigh_op_tnl_2')
// (6, 12, 'neigh_op_lft_2')
// (6, 13, 'neigh_op_bnl_2')

reg n210 = 0;
// (4, 11, 'neigh_op_tnr_3')
// (4, 12, 'neigh_op_rgt_3')
// (4, 13, 'neigh_op_bnr_3')
// (5, 11, 'neigh_op_top_3')
// (5, 12, 'lutff_3/out')
// (5, 12, 'sp4_r_v_b_39')
// (5, 13, 'local_g0_2')
// (5, 13, 'lutff_4/in_0')
// (5, 13, 'neigh_op_bot_3')
// (5, 13, 'sp4_r_v_b_26')
// (5, 14, 'sp4_r_v_b_15')
// (5, 15, 'sp4_r_v_b_2')
// (6, 11, 'neigh_op_tnl_3')
// (6, 11, 'sp4_v_t_39')
// (6, 12, 'neigh_op_lft_3')
// (6, 12, 'sp4_v_b_39')
// (6, 13, 'neigh_op_bnl_3')
// (6, 13, 'sp4_v_b_26')
// (6, 14, 'sp4_v_b_15')
// (6, 15, 'sp4_v_b_2')

reg n211 = 0;
// (4, 11, 'neigh_op_tnr_4')
// (4, 12, 'local_g3_4')
// (4, 12, 'lutff_1/in_0')
// (4, 12, 'neigh_op_rgt_4')
// (4, 13, 'neigh_op_bnr_4')
// (5, 11, 'neigh_op_top_4')
// (5, 12, 'lutff_4/out')
// (5, 13, 'neigh_op_bot_4')
// (6, 11, 'neigh_op_tnl_4')
// (6, 12, 'neigh_op_lft_4')
// (6, 13, 'neigh_op_bnl_4')

reg n212 = 0;
// (4, 11, 'neigh_op_tnr_6')
// (4, 12, 'neigh_op_rgt_6')
// (4, 13, 'neigh_op_bnr_6')
// (5, 11, 'neigh_op_top_6')
// (5, 12, 'lutff_6/out')
// (5, 13, 'local_g1_6')
// (5, 13, 'lutff_3/in_0')
// (5, 13, 'neigh_op_bot_6')
// (6, 11, 'neigh_op_tnl_6')
// (6, 12, 'neigh_op_lft_6')
// (6, 13, 'neigh_op_bnl_6')

reg n213 = 0;
// (4, 11, 'neigh_op_tnr_7')
// (4, 12, 'neigh_op_rgt_7')
// (4, 13, 'neigh_op_bnr_7')
// (5, 11, 'neigh_op_top_7')
// (5, 12, 'local_g1_7')
// (5, 12, 'lutff_6/in_0')
// (5, 12, 'lutff_7/out')
// (5, 13, 'neigh_op_bot_7')
// (6, 11, 'neigh_op_tnl_7')
// (6, 12, 'neigh_op_lft_7')
// (6, 13, 'neigh_op_bnl_7')

reg n214 = 0;
// (4, 11, 'sp12_h_r_1')
// (5, 11, 'sp12_h_r_2')
// (6, 10, 'neigh_op_tnr_7')
// (6, 11, 'neigh_op_rgt_7')
// (6, 11, 'sp12_h_r_5')
// (6, 12, 'neigh_op_bnr_7')
// (7, 10, 'neigh_op_top_7')
// (7, 11, 'lutff_7/out')
// (7, 11, 'sp12_h_r_6')
// (7, 12, 'neigh_op_bot_7')
// (8, 10, 'local_g3_7')
// (8, 10, 'lutff_1/in_1')
// (8, 10, 'neigh_op_tnl_7')
// (8, 11, 'neigh_op_lft_7')
// (8, 11, 'sp12_h_r_9')
// (8, 12, 'neigh_op_bnl_7')
// (9, 11, 'sp12_h_r_10')
// (10, 11, 'sp12_h_r_13')
// (11, 11, 'local_g0_6')
// (11, 11, 'lutff_4/in_0')
// (11, 11, 'sp12_h_r_14')
// (12, 11, 'sp12_h_r_17')
// (13, 11, 'span12_horz_17')

wire n215;
// (4, 12, 'neigh_op_tnr_0')
// (4, 13, 'neigh_op_rgt_0')
// (4, 14, 'neigh_op_bnr_0')
// (5, 12, 'neigh_op_top_0')
// (5, 13, 'lutff_0/out')
// (5, 14, 'neigh_op_bot_0')
// (6, 12, 'local_g3_0')
// (6, 12, 'lutff_0/in_3')
// (6, 12, 'neigh_op_tnl_0')
// (6, 13, 'neigh_op_lft_0')
// (6, 14, 'neigh_op_bnl_0')

wire n216;
// (4, 12, 'neigh_op_tnr_1')
// (4, 13, 'neigh_op_rgt_1')
// (4, 14, 'neigh_op_bnr_1')
// (5, 12, 'neigh_op_top_1')
// (5, 13, 'local_g2_1')
// (5, 13, 'lutff_1/out')
// (5, 13, 'lutff_2/in_3')
// (5, 14, 'neigh_op_bot_1')
// (6, 12, 'neigh_op_tnl_1')
// (6, 13, 'neigh_op_lft_1')
// (6, 14, 'neigh_op_bnl_1')

wire n217;
// (4, 12, 'neigh_op_tnr_2')
// (4, 13, 'neigh_op_rgt_2')
// (4, 14, 'neigh_op_bnr_2')
// (5, 12, 'neigh_op_top_2')
// (5, 13, 'lutff_2/out')
// (5, 14, 'neigh_op_bot_2')
// (6, 12, 'local_g3_2')
// (6, 12, 'lutff_4/in_3')
// (6, 12, 'neigh_op_tnl_2')
// (6, 13, 'neigh_op_lft_2')
// (6, 14, 'neigh_op_bnl_2')

reg n218 = 0;
// (4, 12, 'neigh_op_tnr_3')
// (4, 13, 'neigh_op_rgt_3')
// (4, 14, 'neigh_op_bnr_3')
// (5, 12, 'neigh_op_top_3')
// (5, 13, 'local_g2_3')
// (5, 13, 'lutff_0/in_1')
// (5, 13, 'lutff_3/out')
// (5, 14, 'neigh_op_bot_3')
// (6, 12, 'neigh_op_tnl_3')
// (6, 13, 'local_g0_3')
// (6, 13, 'lutff_6/in_1')
// (6, 13, 'neigh_op_lft_3')
// (6, 14, 'neigh_op_bnl_3')

reg n219 = 0;
// (4, 12, 'neigh_op_tnr_4')
// (4, 13, 'neigh_op_rgt_4')
// (4, 14, 'neigh_op_bnr_4')
// (5, 12, 'neigh_op_top_4')
// (5, 13, 'local_g1_4')
// (5, 13, 'lutff_4/out')
// (5, 13, 'lutff_5/in_0')
// (5, 14, 'neigh_op_bot_4')
// (6, 12, 'neigh_op_tnl_4')
// (6, 13, 'neigh_op_lft_4')
// (6, 14, 'neigh_op_bnl_4')

reg n220 = 0;
// (4, 12, 'neigh_op_tnr_5')
// (4, 12, 'sp4_r_v_b_39')
// (4, 13, 'neigh_op_rgt_5')
// (4, 13, 'sp4_r_v_b_26')
// (4, 14, 'neigh_op_bnr_5')
// (4, 14, 'sp4_r_v_b_15')
// (4, 15, 'sp4_r_v_b_2')
// (5, 11, 'sp4_v_t_39')
// (5, 12, 'neigh_op_top_5')
// (5, 12, 'sp4_v_b_39')
// (5, 13, 'local_g1_5')
// (5, 13, 'lutff_1/in_1')
// (5, 13, 'lutff_5/out')
// (5, 13, 'sp4_v_b_26')
// (5, 14, 'local_g0_7')
// (5, 14, 'lutff_6/in_1')
// (5, 14, 'neigh_op_bot_5')
// (5, 14, 'sp4_v_b_15')
// (5, 15, 'sp4_v_b_2')
// (6, 12, 'neigh_op_tnl_5')
// (6, 13, 'neigh_op_lft_5')
// (6, 14, 'neigh_op_bnl_5')

reg n221 = 0;
// (4, 13, 'neigh_op_tnr_0')
// (4, 14, 'neigh_op_rgt_0')
// (4, 15, 'neigh_op_bnr_0')
// (5, 11, 'sp4_r_v_b_36')
// (5, 12, 'local_g1_1')
// (5, 12, 'lutff_2/in_0')
// (5, 12, 'sp4_r_v_b_25')
// (5, 13, 'local_g0_0')
// (5, 13, 'lutff_2/in_0')
// (5, 13, 'neigh_op_top_0')
// (5, 13, 'sp4_r_v_b_12')
// (5, 14, 'local_g0_0')
// (5, 14, 'lutff_0/out')
// (5, 14, 'lutff_4/in_0')
// (5, 14, 'lutff_6/in_0')
// (5, 14, 'sp4_r_v_b_1')
// (5, 15, 'neigh_op_bot_0')
// (6, 10, 'sp4_v_t_36')
// (6, 11, 'sp4_v_b_36')
// (6, 12, 'sp4_v_b_25')
// (6, 13, 'neigh_op_tnl_0')
// (6, 13, 'sp4_v_b_12')
// (6, 14, 'neigh_op_lft_0')
// (6, 14, 'sp4_v_b_1')
// (6, 15, 'neigh_op_bnl_0')

reg n222 = 0;
// (4, 13, 'neigh_op_tnr_1')
// (4, 14, 'neigh_op_rgt_1')
// (4, 15, 'neigh_op_bnr_1')
// (5, 13, 'local_g0_1')
// (5, 13, 'lutff_1/in_0')
// (5, 13, 'neigh_op_top_1')
// (5, 14, 'local_g0_1')
// (5, 14, 'lutff_1/out')
// (5, 14, 'lutff_4/in_1')
// (5, 15, 'neigh_op_bot_1')
// (6, 13, 'neigh_op_tnl_1')
// (6, 14, 'neigh_op_lft_1')
// (6, 15, 'neigh_op_bnl_1')

reg n223 = 0;
// (4, 13, 'neigh_op_tnr_2')
// (4, 14, 'neigh_op_rgt_2')
// (4, 15, 'neigh_op_bnr_2')
// (5, 13, 'neigh_op_top_2')
// (5, 14, 'local_g1_2')
// (5, 14, 'lutff_1/in_0')
// (5, 14, 'lutff_2/out')
// (5, 15, 'neigh_op_bot_2')
// (6, 13, 'neigh_op_tnl_2')
// (6, 14, 'neigh_op_lft_2')
// (6, 15, 'neigh_op_bnl_2')

reg n224 = 0;
// (4, 13, 'neigh_op_tnr_6')
// (4, 14, 'neigh_op_rgt_6')
// (4, 15, 'neigh_op_bnr_6')
// (5, 13, 'neigh_op_top_6')
// (5, 14, 'local_g1_6')
// (5, 14, 'lutff_6/out')
// (5, 14, 'lutff_7/in_0')
// (5, 15, 'neigh_op_bot_6')
// (6, 13, 'neigh_op_tnl_6')
// (6, 14, 'neigh_op_lft_6')
// (6, 15, 'neigh_op_bnl_6')

reg n225 = 0;
// (4, 13, 'neigh_op_tnr_7')
// (4, 14, 'neigh_op_rgt_7')
// (4, 15, 'neigh_op_bnr_7')
// (5, 13, 'neigh_op_top_7')
// (5, 14, 'local_g1_7')
// (5, 14, 'lutff_2/in_0')
// (5, 14, 'lutff_7/out')
// (5, 15, 'neigh_op_bot_7')
// (6, 13, 'neigh_op_tnl_7')
// (6, 14, 'neigh_op_lft_7')
// (6, 15, 'neigh_op_bnl_7')

wire n226;
// (5, 1, 'neigh_op_tnr_7')
// (5, 2, 'neigh_op_rgt_7')
// (5, 3, 'neigh_op_bnr_7')
// (6, 1, 'neigh_op_top_7')
// (6, 2, 'lutff_7/out')
// (6, 3, 'neigh_op_bot_7')
// (7, 1, 'neigh_op_tnl_7')
// (7, 2, 'local_g1_7')
// (7, 2, 'lutff_1/in_3')
// (7, 2, 'neigh_op_lft_7')
// (7, 3, 'neigh_op_bnl_7')

wire n227;
// (5, 1, 'sp4_r_v_b_24')
// (5, 2, 'neigh_op_tnr_0')
// (5, 2, 'sp4_r_v_b_13')
// (5, 3, 'neigh_op_rgt_0')
// (5, 3, 'sp4_r_v_b_0')
// (5, 4, 'neigh_op_bnr_0')
// (6, 0, 'span4_vert_24')
// (6, 1, 'sp4_r_v_b_25')
// (6, 1, 'sp4_v_b_24')
// (6, 2, 'local_g1_5')
// (6, 2, 'lutff_7/in_3')
// (6, 2, 'neigh_op_top_0')
// (6, 2, 'sp4_r_v_b_12')
// (6, 2, 'sp4_v_b_13')
// (6, 3, 'lutff_0/out')
// (6, 3, 'sp4_r_v_b_1')
// (6, 3, 'sp4_v_b_0')
// (6, 4, 'neigh_op_bot_0')
// (7, 0, 'span4_vert_25')
// (7, 1, 'sp4_v_b_25')
// (7, 2, 'local_g0_4')
// (7, 2, 'lutff_0/in_2')
// (7, 2, 'lutff_6/in_2')
// (7, 2, 'neigh_op_tnl_0')
// (7, 2, 'sp4_v_b_12')
// (7, 3, 'local_g1_0')
// (7, 3, 'lutff_0/in_3')
// (7, 3, 'neigh_op_lft_0')
// (7, 3, 'sp4_h_r_7')
// (7, 3, 'sp4_v_b_1')
// (7, 4, 'neigh_op_bnl_0')
// (8, 3, 'local_g0_2')
// (8, 3, 'lutff_4/in_2')
// (8, 3, 'sp4_h_r_18')
// (9, 3, 'sp4_h_r_31')
// (10, 3, 'sp4_h_r_42')
// (11, 3, 'sp4_h_l_42')

reg n228 = 0;
// (5, 1, 'sp4_r_v_b_43')
// (5, 2, 'sp4_r_v_b_30')
// (5, 3, 'sp4_r_v_b_19')
// (5, 4, 'sp4_r_v_b_6')
// (6, 0, 'span4_vert_43')
// (6, 1, 'sp4_v_b_43')
// (6, 2, 'sp4_v_b_30')
// (6, 3, 'local_g0_3')
// (6, 3, 'lutff_7/in_0')
// (6, 3, 'sp4_v_b_19')
// (6, 4, 'sp4_h_r_6')
// (6, 4, 'sp4_v_b_6')
// (6, 10, 'sp4_h_r_9')
// (7, 4, 'sp4_h_r_19')
// (7, 10, 'local_g0_4')
// (7, 10, 'local_g1_4')
// (7, 10, 'lutff_4/in_2')
// (7, 10, 'lutff_5/in_2')
// (7, 10, 'sp4_h_r_20')
// (8, 3, 'neigh_op_tnr_0')
// (8, 4, 'neigh_op_rgt_0')
// (8, 4, 'sp4_h_r_30')
// (8, 5, 'neigh_op_bnr_0')
// (8, 10, 'sp4_h_r_33')
// (9, 1, 'sp4_r_v_b_36')
// (9, 2, 'sp4_r_v_b_25')
// (9, 3, 'neigh_op_top_0')
// (9, 3, 'sp4_r_v_b_12')
// (9, 3, 'sp4_r_v_b_44')
// (9, 4, 'lutff_0/out')
// (9, 4, 'sp4_h_r_43')
// (9, 4, 'sp4_r_v_b_1')
// (9, 4, 'sp4_r_v_b_33')
// (9, 5, 'neigh_op_bot_0')
// (9, 5, 'sp4_r_v_b_20')
// (9, 6, 'sp4_r_v_b_9')
// (9, 7, 'sp4_r_v_b_44')
// (9, 8, 'sp4_r_v_b_33')
// (9, 9, 'sp4_r_v_b_20')
// (9, 10, 'sp4_h_r_44')
// (9, 10, 'sp4_r_v_b_9')
// (10, 0, 'span4_vert_36')
// (10, 1, 'sp4_v_b_36')
// (10, 2, 'sp4_v_b_25')
// (10, 2, 'sp4_v_t_44')
// (10, 3, 'neigh_op_tnl_0')
// (10, 3, 'sp4_v_b_12')
// (10, 3, 'sp4_v_b_44')
// (10, 4, 'neigh_op_lft_0')
// (10, 4, 'sp4_h_l_43')
// (10, 4, 'sp4_v_b_1')
// (10, 4, 'sp4_v_b_33')
// (10, 5, 'neigh_op_bnl_0')
// (10, 5, 'sp4_v_b_20')
// (10, 6, 'sp4_v_b_9')
// (10, 6, 'sp4_v_t_44')
// (10, 7, 'sp4_v_b_44')
// (10, 8, 'sp4_v_b_33')
// (10, 9, 'sp4_v_b_20')
// (10, 10, 'sp4_h_l_44')
// (10, 10, 'sp4_h_r_0')
// (10, 10, 'sp4_v_b_9')
// (11, 10, 'sp4_h_r_13')
// (12, 10, 'local_g2_0')
// (12, 10, 'lutff_0/in_0')
// (12, 10, 'sp4_h_r_24')
// (13, 10, 'span4_horz_24')

wire n229;
// (5, 2, 'neigh_op_tnr_2')
// (5, 3, 'neigh_op_rgt_2')
// (5, 4, 'neigh_op_bnr_2')
// (6, 2, 'neigh_op_top_2')
// (6, 3, 'local_g0_2')
// (6, 3, 'lutff_0/in_2')
// (6, 3, 'lutff_2/out')
// (6, 3, 'sp4_r_v_b_37')
// (6, 4, 'local_g0_0')
// (6, 4, 'local_g1_2')
// (6, 4, 'lutff_1/in_0')
// (6, 4, 'lutff_5/in_1')
// (6, 4, 'neigh_op_bot_2')
// (6, 4, 'sp4_r_v_b_24')
// (6, 5, 'sp4_r_v_b_13')
// (6, 6, 'sp4_r_v_b_0')
// (7, 2, 'neigh_op_tnl_2')
// (7, 2, 'sp4_v_t_37')
// (7, 3, 'neigh_op_lft_2')
// (7, 3, 'sp4_v_b_37')
// (7, 4, 'neigh_op_bnl_2')
// (7, 4, 'sp4_v_b_24')
// (7, 5, 'sp4_v_b_13')
// (7, 6, 'sp4_v_b_0')

wire n230;
// (5, 2, 'neigh_op_tnr_4')
// (5, 2, 'sp4_r_v_b_37')
// (5, 3, 'neigh_op_rgt_4')
// (5, 3, 'sp4_r_v_b_24')
// (5, 4, 'neigh_op_bnr_4')
// (5, 4, 'sp4_r_v_b_13')
// (5, 5, 'sp4_r_v_b_0')
// (6, 1, 'sp4_v_t_37')
// (6, 2, 'neigh_op_top_4')
// (6, 2, 'sp4_v_b_37')
// (6, 3, 'lutff_4/out')
// (6, 3, 'sp4_v_b_24')
// (6, 4, 'local_g0_5')
// (6, 4, 'lutff_1/in_2')
// (6, 4, 'lutff_6/in_3')
// (6, 4, 'neigh_op_bot_4')
// (6, 4, 'sp4_v_b_13')
// (6, 5, 'sp4_v_b_0')
// (7, 2, 'neigh_op_tnl_4')
// (7, 3, 'neigh_op_lft_4')
// (7, 4, 'neigh_op_bnl_4')

reg n231 = 0;
// (5, 2, 'neigh_op_tnr_7')
// (5, 3, 'neigh_op_rgt_7')
// (5, 4, 'neigh_op_bnr_7')
// (6, 2, 'neigh_op_top_7')
// (6, 3, 'local_g2_7')
// (6, 3, 'lutff_4/in_3')
// (6, 3, 'lutff_7/out')
// (6, 4, 'neigh_op_bot_7')
// (7, 2, 'neigh_op_tnl_7')
// (7, 3, 'neigh_op_lft_7')
// (7, 4, 'neigh_op_bnl_7')

wire n232;
// (5, 3, 'neigh_op_tnr_1')
// (5, 4, 'neigh_op_rgt_1')
// (5, 5, 'neigh_op_bnr_1')
// (6, 3, 'neigh_op_top_1')
// (6, 4, 'local_g1_1')
// (6, 4, 'lutff_0/in_2')
// (6, 4, 'lutff_1/out')
// (6, 4, 'lutff_2/in_2')
// (6, 5, 'local_g1_1')
// (6, 5, 'lutff_7/in_3')
// (6, 5, 'neigh_op_bot_1')
// (7, 3, 'neigh_op_tnl_1')
// (7, 4, 'neigh_op_lft_1')
// (7, 5, 'neigh_op_bnl_1')

wire n233;
// (5, 3, 'neigh_op_tnr_2')
// (5, 4, 'neigh_op_rgt_2')
// (5, 5, 'neigh_op_bnr_2')
// (6, 3, 'neigh_op_top_2')
// (6, 4, 'lutff_2/out')
// (6, 4, 'sp4_h_r_4')
// (6, 5, 'neigh_op_bot_2')
// (7, 3, 'local_g2_2')
// (7, 3, 'lutff_5/in_3')
// (7, 3, 'lutff_7/in_3')
// (7, 3, 'neigh_op_tnl_2')
// (7, 4, 'local_g1_1')
// (7, 4, 'lutff_7/in_3')
// (7, 4, 'neigh_op_lft_2')
// (7, 4, 'sp4_h_r_17')
// (7, 5, 'neigh_op_bnl_2')
// (8, 4, 'local_g2_4')
// (8, 4, 'lutff_2/in_2')
// (8, 4, 'sp4_h_r_28')
// (9, 4, 'sp4_h_r_41')
// (10, 4, 'sp4_h_l_41')

wire n234;
// (5, 3, 'neigh_op_tnr_3')
// (5, 4, 'neigh_op_rgt_3')
// (5, 5, 'neigh_op_bnr_3')
// (6, 3, 'neigh_op_top_3')
// (6, 4, 'local_g1_3')
// (6, 4, 'lutff_1/in_1')
// (6, 4, 'lutff_3/out')
// (6, 4, 'lutff_6/in_2')
// (6, 5, 'neigh_op_bot_3')
// (7, 3, 'neigh_op_tnl_3')
// (7, 4, 'neigh_op_lft_3')
// (7, 5, 'neigh_op_bnl_3')

wire n235;
// (5, 3, 'neigh_op_tnr_4')
// (5, 4, 'neigh_op_rgt_4')
// (5, 5, 'neigh_op_bnr_4')
// (6, 3, 'neigh_op_top_4')
// (6, 4, 'lutff_4/out')
// (6, 4, 'sp4_h_r_8')
// (6, 4, 'sp4_r_v_b_41')
// (6, 5, 'neigh_op_bot_4')
// (6, 5, 'sp4_r_v_b_28')
// (6, 6, 'sp4_r_v_b_17')
// (6, 7, 'sp4_r_v_b_4')
// (7, 3, 'local_g2_4')
// (7, 3, 'lutff_2/in_2')
// (7, 3, 'lutff_7/in_1')
// (7, 3, 'neigh_op_tnl_4')
// (7, 3, 'sp4_h_r_4')
// (7, 3, 'sp4_h_r_9')
// (7, 3, 'sp4_v_t_41')
// (7, 4, 'neigh_op_lft_4')
// (7, 4, 'sp4_h_r_21')
// (7, 4, 'sp4_v_b_41')
// (7, 5, 'neigh_op_bnl_4')
// (7, 5, 'sp4_v_b_28')
// (7, 6, 'sp4_v_b_17')
// (7, 7, 'sp4_v_b_4')
// (8, 3, 'local_g1_1')
// (8, 3, 'local_g1_4')
// (8, 3, 'lutff_1/in_3')
// (8, 3, 'lutff_7/in_2')
// (8, 3, 'sp4_h_r_17')
// (8, 3, 'sp4_h_r_20')
// (8, 4, 'local_g3_0')
// (8, 4, 'lutff_7/in_2')
// (8, 4, 'sp4_h_r_32')
// (9, 3, 'sp4_h_r_28')
// (9, 3, 'sp4_h_r_33')
// (9, 4, 'sp4_h_r_45')
// (10, 3, 'sp4_h_r_41')
// (10, 3, 'sp4_h_r_44')
// (10, 4, 'sp4_h_l_45')
// (11, 3, 'sp4_h_l_41')
// (11, 3, 'sp4_h_l_44')

wire n236;
// (5, 3, 'neigh_op_tnr_5')
// (5, 4, 'neigh_op_rgt_5')
// (5, 5, 'neigh_op_bnr_5')
// (6, 3, 'neigh_op_top_5')
// (6, 4, 'lutff_5/out')
// (6, 5, 'neigh_op_bot_5')
// (7, 3, 'neigh_op_tnl_5')
// (7, 4, 'local_g0_5')
// (7, 4, 'local_g1_5')
// (7, 4, 'lutff_0/in_1')
// (7, 4, 'lutff_2/in_2')
// (7, 4, 'lutff_4/in_2')
// (7, 4, 'lutff_6/in_1')
// (7, 4, 'neigh_op_lft_5')
// (7, 5, 'neigh_op_bnl_5')

wire n237;
// (5, 3, 'neigh_op_tnr_7')
// (5, 4, 'neigh_op_rgt_7')
// (5, 5, 'neigh_op_bnr_7')
// (6, 3, 'neigh_op_top_7')
// (6, 4, 'local_g0_7')
// (6, 4, 'local_g1_7')
// (6, 4, 'lutff_0/in_1')
// (6, 4, 'lutff_2/in_0')
// (6, 4, 'lutff_4/in_1')
// (6, 4, 'lutff_7/out')
// (6, 5, 'neigh_op_bot_7')
// (7, 3, 'neigh_op_tnl_7')
// (7, 4, 'neigh_op_lft_7')
// (7, 5, 'neigh_op_bnl_7')

reg n238 = 0;
// (5, 3, 'sp4_h_r_2')
// (6, 3, 'local_g0_7')
// (6, 3, 'lutff_2/in_3')
// (6, 3, 'sp4_h_r_15')
// (7, 3, 'sp4_h_r_26')
// (8, 2, 'neigh_op_tnr_3')
// (8, 3, 'neigh_op_rgt_3')
// (8, 3, 'sp4_h_r_39')
// (8, 4, 'neigh_op_bnr_3')
// (9, 2, 'neigh_op_top_3')
// (9, 3, 'local_g0_3')
// (9, 3, 'lutff_3/out')
// (9, 3, 'lutff_7/in_0')
// (9, 3, 'sp4_h_l_39')
// (9, 3, 'sp4_h_r_6')
// (9, 4, 'neigh_op_bot_3')
// (10, 2, 'neigh_op_tnl_3')
// (10, 3, 'neigh_op_lft_3')
// (10, 3, 'sp4_h_r_19')
// (10, 4, 'neigh_op_bnl_3')
// (11, 3, 'sp4_h_r_30')
// (12, 3, 'sp4_h_r_43')
// (13, 3, 'span4_horz_43')

wire n239;
// (5, 3, 'sp4_r_v_b_38')
// (5, 4, 'neigh_op_tnr_7')
// (5, 4, 'sp4_r_v_b_27')
// (5, 5, 'neigh_op_rgt_7')
// (5, 5, 'sp4_r_v_b_14')
// (5, 6, 'neigh_op_bnr_7')
// (5, 6, 'sp4_r_v_b_3')
// (6, 1, 'sp4_r_v_b_31')
// (6, 2, 'sp4_r_v_b_18')
// (6, 2, 'sp4_v_t_38')
// (6, 3, 'local_g3_6')
// (6, 3, 'lutff_6/in_3')
// (6, 3, 'sp4_r_v_b_7')
// (6, 3, 'sp4_v_b_38')
// (6, 4, 'neigh_op_top_7')
// (6, 4, 'sp4_r_v_b_42')
// (6, 4, 'sp4_v_b_27')
// (6, 5, 'lutff_7/out')
// (6, 5, 'sp4_r_v_b_31')
// (6, 5, 'sp4_v_b_14')
// (6, 6, 'neigh_op_bot_7')
// (6, 6, 'sp4_r_v_b_18')
// (6, 6, 'sp4_v_b_3')
// (6, 7, 'sp4_r_v_b_7')
// (7, 0, 'span4_vert_31')
// (7, 1, 'sp4_v_b_31')
// (7, 2, 'sp4_v_b_18')
// (7, 3, 'local_g0_7')
// (7, 3, 'lutff_7/in_2')
// (7, 3, 'sp4_v_b_7')
// (7, 3, 'sp4_v_t_42')
// (7, 4, 'local_g3_7')
// (7, 4, 'lutff_5/in_3')
// (7, 4, 'neigh_op_tnl_7')
// (7, 4, 'sp4_v_b_42')
// (7, 5, 'neigh_op_lft_7')
// (7, 5, 'sp4_v_b_31')
// (7, 6, 'neigh_op_bnl_7')
// (7, 6, 'sp4_v_b_18')
// (7, 7, 'sp4_v_b_7')

reg n240 = 0;
// (5, 3, 'sp4_r_v_b_39')
// (5, 4, 'sp4_r_v_b_26')
// (5, 5, 'neigh_op_tnr_1')
// (5, 5, 'sp4_r_v_b_15')
// (5, 6, 'neigh_op_rgt_1')
// (5, 6, 'sp4_r_v_b_2')
// (5, 7, 'neigh_op_bnr_1')
// (6, 2, 'sp4_v_t_39')
// (6, 3, 'sp4_v_b_39')
// (6, 4, 'sp4_v_b_26')
// (6, 5, 'local_g0_7')
// (6, 5, 'lutff_2/in_3')
// (6, 5, 'neigh_op_top_1')
// (6, 5, 'sp4_v_b_15')
// (6, 6, 'lutff_1/out')
// (6, 6, 'sp4_v_b_2')
// (6, 7, 'neigh_op_bot_1')
// (7, 5, 'neigh_op_tnl_1')
// (7, 6, 'neigh_op_lft_1')
// (7, 7, 'neigh_op_bnl_1')

wire n241;
// (5, 4, 'neigh_op_tnr_0')
// (5, 5, 'neigh_op_rgt_0')
// (5, 6, 'neigh_op_bnr_0')
// (6, 4, 'neigh_op_top_0')
// (6, 5, 'local_g0_0')
// (6, 5, 'lutff_0/out')
// (6, 5, 'lutff_5/in_1')
// (6, 5, 'lutff_7/in_1')
// (6, 6, 'neigh_op_bot_0')
// (7, 4, 'neigh_op_tnl_0')
// (7, 5, 'neigh_op_lft_0')
// (7, 6, 'neigh_op_bnl_0')

wire n242;
// (5, 4, 'neigh_op_tnr_1')
// (5, 5, 'neigh_op_rgt_1')
// (5, 6, 'neigh_op_bnr_1')
// (6, 4, 'neigh_op_top_1')
// (6, 5, 'local_g0_1')
// (6, 5, 'lutff_1/out')
// (6, 5, 'lutff_5/in_2')
// (6, 5, 'lutff_7/in_2')
// (6, 6, 'neigh_op_bot_1')
// (7, 4, 'neigh_op_tnl_1')
// (7, 5, 'neigh_op_lft_1')
// (7, 6, 'neigh_op_bnl_1')

wire n243;
// (5, 4, 'neigh_op_tnr_2')
// (5, 5, 'neigh_op_rgt_2')
// (5, 6, 'neigh_op_bnr_2')
// (6, 4, 'local_g0_2')
// (6, 4, 'lutff_5/in_3')
// (6, 4, 'lutff_7/in_3')
// (6, 4, 'neigh_op_top_2')
// (6, 5, 'lutff_2/out')
// (6, 6, 'neigh_op_bot_2')
// (7, 4, 'neigh_op_tnl_2')
// (7, 5, 'neigh_op_lft_2')
// (7, 6, 'neigh_op_bnl_2')

wire n244;
// (5, 4, 'neigh_op_tnr_3')
// (5, 5, 'neigh_op_rgt_3')
// (5, 6, 'neigh_op_bnr_3')
// (6, 4, 'neigh_op_top_3')
// (6, 5, 'lutff_3/out')
// (6, 6, 'neigh_op_bot_3')
// (7, 4, 'neigh_op_tnl_3')
// (7, 5, 'local_g1_3')
// (7, 5, 'lutff_1/in_3')
// (7, 5, 'neigh_op_lft_3')
// (7, 6, 'neigh_op_bnl_3')

wire n245;
// (5, 4, 'neigh_op_tnr_4')
// (5, 5, 'neigh_op_rgt_4')
// (5, 6, 'neigh_op_bnr_4')
// (6, 4, 'neigh_op_top_4')
// (6, 5, 'local_g0_4')
// (6, 5, 'local_g1_4')
// (6, 5, 'lutff_4/out')
// (6, 5, 'lutff_5/in_3')
// (6, 5, 'lutff_6/in_3')
// (6, 6, 'neigh_op_bot_4')
// (7, 4, 'neigh_op_tnl_4')
// (7, 5, 'neigh_op_lft_4')
// (7, 6, 'neigh_op_bnl_4')

wire n246;
// (5, 4, 'neigh_op_tnr_5')
// (5, 5, 'neigh_op_rgt_5')
// (5, 6, 'neigh_op_bnr_5')
// (6, 0, 'span12_vert_18')
// (6, 1, 'sp12_v_b_18')
// (6, 2, 'sp12_v_b_17')
// (6, 3, 'sp12_v_b_14')
// (6, 4, 'local_g2_5')
// (6, 4, 'lutff_0/in_3')
// (6, 4, 'lutff_4/in_3')
// (6, 4, 'neigh_op_top_5')
// (6, 4, 'sp12_v_b_13')
// (6, 5, 'lutff_5/out')
// (6, 5, 'sp12_v_b_10')
// (6, 6, 'neigh_op_bot_5')
// (6, 6, 'sp12_v_b_9')
// (6, 7, 'sp12_v_b_6')
// (6, 8, 'sp12_v_b_5')
// (6, 9, 'sp12_v_b_2')
// (6, 10, 'sp12_v_b_1')
// (7, 4, 'neigh_op_tnl_5')
// (7, 5, 'neigh_op_lft_5')
// (7, 6, 'neigh_op_bnl_5')

wire n247;
// (5, 4, 'neigh_op_tnr_6')
// (5, 5, 'neigh_op_rgt_6')
// (5, 6, 'neigh_op_bnr_6')
// (6, 4, 'local_g1_6')
// (6, 4, 'lutff_2/in_3')
// (6, 4, 'neigh_op_top_6')
// (6, 5, 'lutff_6/out')
// (6, 6, 'neigh_op_bot_6')
// (7, 4, 'neigh_op_tnl_6')
// (7, 5, 'neigh_op_lft_6')
// (7, 6, 'neigh_op_bnl_6')

wire n248;
// (5, 4, 'sp4_h_r_6')
// (6, 3, 'neigh_op_tnr_7')
// (6, 4, 'neigh_op_rgt_7')
// (6, 4, 'sp4_h_r_19')
// (6, 5, 'neigh_op_bnr_7')
// (7, 3, 'local_g1_7')
// (7, 3, 'lutff_0/in_0')
// (7, 3, 'lutff_6/in_0')
// (7, 3, 'neigh_op_top_7')
// (7, 4, 'lutff_7/out')
// (7, 4, 'sp4_h_r_30')
// (7, 5, 'neigh_op_bot_7')
// (8, 3, 'local_g2_7')
// (8, 3, 'lutff_1/in_0')
// (8, 3, 'neigh_op_tnl_7')
// (8, 4, 'local_g2_3')
// (8, 4, 'local_g3_3')
// (8, 4, 'lutff_4/in_3')
// (8, 4, 'lutff_5/in_3')
// (8, 4, 'neigh_op_lft_7')
// (8, 4, 'sp4_h_r_43')
// (8, 5, 'neigh_op_bnl_7')
// (9, 4, 'sp4_h_l_43')

wire n249;
// (5, 4, 'sp4_h_r_8')
// (6, 4, 'sp4_h_r_21')
// (7, 1, 'neigh_op_tnr_5')
// (7, 2, 'neigh_op_rgt_5')
// (7, 3, 'neigh_op_bnr_5')
// (7, 4, 'sp4_h_r_32')
// (8, 1, 'neigh_op_top_5')
// (8, 1, 'sp4_r_v_b_38')
// (8, 2, 'lutff_5/out')
// (8, 2, 'sp4_r_v_b_27')
// (8, 3, 'local_g0_5')
// (8, 3, 'lutff_7/in_0')
// (8, 3, 'neigh_op_bot_5')
// (8, 3, 'sp4_r_v_b_14')
// (8, 4, 'local_g1_3')
// (8, 4, 'local_g2_5')
// (8, 4, 'lutff_4/in_0')
// (8, 4, 'lutff_5/in_0')
// (8, 4, 'lutff_7/in_0')
// (8, 4, 'sp4_h_r_45')
// (8, 4, 'sp4_r_v_b_3')
// (9, 0, 'span4_vert_38')
// (9, 1, 'neigh_op_tnl_5')
// (9, 1, 'sp4_v_b_38')
// (9, 2, 'neigh_op_lft_5')
// (9, 2, 'sp4_v_b_27')
// (9, 3, 'neigh_op_bnl_5')
// (9, 3, 'sp4_v_b_14')
// (9, 4, 'sp4_h_l_45')
// (9, 4, 'sp4_v_b_3')

reg n250 = 0;
// (5, 5, 'local_g3_5')
// (5, 5, 'lutff_1/in_3')
// (5, 5, 'neigh_op_tnr_5')
// (5, 6, 'neigh_op_rgt_5')
// (5, 7, 'neigh_op_bnr_5')
// (6, 5, 'neigh_op_top_5')
// (6, 6, 'lutff_5/out')
// (6, 7, 'neigh_op_bot_5')
// (7, 5, 'neigh_op_tnl_5')
// (7, 6, 'neigh_op_lft_5')
// (7, 7, 'neigh_op_bnl_5')

reg n251 = 0;
// (5, 5, 'neigh_op_tnr_2')
// (5, 6, 'neigh_op_rgt_2')
// (5, 7, 'neigh_op_bnr_2')
// (6, 5, 'local_g1_2')
// (6, 5, 'lutff_4/in_3')
// (6, 5, 'neigh_op_top_2')
// (6, 6, 'lutff_2/out')
// (6, 7, 'neigh_op_bot_2')
// (7, 5, 'neigh_op_tnl_2')
// (7, 6, 'neigh_op_lft_2')
// (7, 7, 'neigh_op_bnl_2')

reg n252 = 0;
// (5, 5, 'neigh_op_tnr_6')
// (5, 6, 'neigh_op_rgt_6')
// (5, 7, 'neigh_op_bnr_6')
// (6, 5, 'local_g0_6')
// (6, 5, 'lutff_1/in_3')
// (6, 5, 'neigh_op_top_6')
// (6, 6, 'lutff_6/out')
// (6, 7, 'neigh_op_bot_6')
// (7, 5, 'neigh_op_tnl_6')
// (7, 6, 'neigh_op_lft_6')
// (7, 7, 'neigh_op_bnl_6')

wire n253;
// (5, 5, 'sp4_h_r_9')
// (6, 5, 'sp4_h_r_20')
// (7, 2, 'neigh_op_tnr_0')
// (7, 3, 'neigh_op_rgt_0')
// (7, 4, 'neigh_op_bnr_0')
// (7, 5, 'sp4_h_r_33')
// (8, 2, 'neigh_op_top_0')
// (8, 2, 'sp4_r_v_b_44')
// (8, 3, 'lutff_0/out')
// (8, 3, 'sp4_r_v_b_33')
// (8, 4, 'neigh_op_bot_0')
// (8, 4, 'sp4_r_v_b_20')
// (8, 5, 'local_g2_1')
// (8, 5, 'local_g2_4')
// (8, 5, 'lutff_2/in_3')
// (8, 5, 'lutff_3/in_3')
// (8, 5, 'lutff_5/in_2')
// (8, 5, 'sp4_h_r_44')
// (8, 5, 'sp4_r_v_b_9')
// (9, 1, 'sp4_v_t_44')
// (9, 2, 'neigh_op_tnl_0')
// (9, 2, 'sp4_v_b_44')
// (9, 3, 'neigh_op_lft_0')
// (9, 3, 'sp4_v_b_33')
// (9, 4, 'neigh_op_bnl_0')
// (9, 4, 'sp4_v_b_20')
// (9, 5, 'sp4_h_l_44')
// (9, 5, 'sp4_v_b_9')

wire n254;
// (5, 5, 'sp4_r_v_b_47')
// (5, 6, 'sp4_r_v_b_34')
// (5, 7, 'neigh_op_tnr_5')
// (5, 7, 'sp4_r_v_b_23')
// (5, 8, 'neigh_op_rgt_5')
// (5, 8, 'sp4_r_v_b_10')
// (5, 9, 'neigh_op_bnr_5')
// (6, 4, 'sp4_v_t_47')
// (6, 5, 'sp4_v_b_47')
// (6, 6, 'sp4_v_b_34')
// (6, 7, 'local_g0_5')
// (6, 7, 'local_g1_7')
// (6, 7, 'lutff_3/in_2')
// (6, 7, 'lutff_7/in_3')
// (6, 7, 'neigh_op_top_5')
// (6, 7, 'sp4_v_b_23')
// (6, 8, 'lutff_5/out')
// (6, 8, 'sp4_r_v_b_43')
// (6, 8, 'sp4_v_b_10')
// (6, 9, 'neigh_op_bot_5')
// (6, 9, 'sp4_r_v_b_30')
// (6, 10, 'sp4_r_v_b_19')
// (6, 11, 'sp4_r_v_b_6')
// (7, 7, 'local_g2_5')
// (7, 7, 'local_g3_5')
// (7, 7, 'lutff_0/in_3')
// (7, 7, 'lutff_6/in_2')
// (7, 7, 'neigh_op_tnl_5')
// (7, 7, 'sp4_h_r_6')
// (7, 7, 'sp4_v_t_43')
// (7, 8, 'local_g1_5')
// (7, 8, 'lutff_5/in_1')
// (7, 8, 'neigh_op_lft_5')
// (7, 8, 'sp4_v_b_43')
// (7, 9, 'neigh_op_bnl_5')
// (7, 9, 'sp4_v_b_30')
// (7, 10, 'sp4_v_b_19')
// (7, 11, 'sp4_v_b_6')
// (8, 7, 'local_g1_3')
// (8, 7, 'lutff_0/in_2')
// (8, 7, 'lutff_3/in_1')
// (8, 7, 'lutff_5/in_1')
// (8, 7, 'sp4_h_r_19')
// (9, 7, 'sp4_h_r_30')
// (10, 7, 'sp4_h_r_43')
// (11, 7, 'sp4_h_l_43')

wire n255;
// (5, 6, 'neigh_op_tnr_2')
// (5, 7, 'neigh_op_rgt_2')
// (5, 7, 'sp4_h_r_9')
// (5, 8, 'neigh_op_bnr_2')
// (6, 5, 'sp4_r_v_b_45')
// (6, 6, 'neigh_op_top_2')
// (6, 6, 'sp4_r_v_b_32')
// (6, 7, 'lutff_2/out')
// (6, 7, 'sp4_h_r_20')
// (6, 7, 'sp4_r_v_b_21')
// (6, 7, 'sp4_r_v_b_37')
// (6, 8, 'neigh_op_bot_2')
// (6, 8, 'sp4_r_v_b_24')
// (6, 8, 'sp4_r_v_b_8')
// (6, 9, 'sp4_r_v_b_13')
// (6, 10, 'sp4_r_v_b_0')
// (7, 4, 'sp4_v_t_45')
// (7, 5, 'sp4_v_b_45')
// (7, 6, 'neigh_op_tnl_2')
// (7, 6, 'sp4_h_r_5')
// (7, 6, 'sp4_v_b_32')
// (7, 6, 'sp4_v_t_37')
// (7, 7, 'neigh_op_lft_2')
// (7, 7, 'sp4_h_r_33')
// (7, 7, 'sp4_v_b_21')
// (7, 7, 'sp4_v_b_37')
// (7, 8, 'local_g0_0')
// (7, 8, 'local_g3_2')
// (7, 8, 'lutff_0/in_0')
// (7, 8, 'lutff_6/in_2')
// (7, 8, 'lutff_7/in_0')
// (7, 8, 'neigh_op_bnl_2')
// (7, 8, 'sp4_v_b_24')
// (7, 8, 'sp4_v_b_8')
// (7, 9, 'sp4_v_b_13')
// (7, 10, 'sp4_v_b_0')
// (8, 4, 'sp4_r_v_b_44')
// (8, 5, 'sp4_r_v_b_33')
// (8, 6, 'local_g0_0')
// (8, 6, 'local_g3_4')
// (8, 6, 'lutff_2/in_2')
// (8, 6, 'lutff_4/in_1')
// (8, 6, 'lutff_5/in_0')
// (8, 6, 'lutff_6/in_1')
// (8, 6, 'sp4_h_r_16')
// (8, 6, 'sp4_r_v_b_20')
// (8, 7, 'local_g3_4')
// (8, 7, 'lutff_1/in_2')
// (8, 7, 'sp4_h_r_44')
// (8, 7, 'sp4_r_v_b_9')
// (9, 3, 'sp4_v_t_44')
// (9, 4, 'sp4_v_b_44')
// (9, 5, 'sp4_v_b_33')
// (9, 6, 'sp4_h_r_29')
// (9, 6, 'sp4_v_b_20')
// (9, 7, 'sp4_h_l_44')
// (9, 7, 'sp4_v_b_9')
// (10, 6, 'sp4_h_r_40')
// (11, 6, 'sp4_h_l_40')

wire n256;
// (5, 6, 'neigh_op_tnr_3')
// (5, 7, 'neigh_op_rgt_3')
// (5, 8, 'neigh_op_bnr_3')
// (6, 6, 'neigh_op_top_3')
// (6, 6, 'sp12_h_r_1')
// (6, 6, 'sp12_v_t_22')
// (6, 7, 'local_g0_3')
// (6, 7, 'lutff_2/in_1')
// (6, 7, 'lutff_3/out')
// (6, 7, 'sp12_v_b_22')
// (6, 8, 'neigh_op_bot_3')
// (6, 8, 'sp12_v_b_21')
// (6, 9, 'sp12_v_b_18')
// (6, 10, 'sp12_v_b_17')
// (6, 11, 'sp12_v_b_14')
// (6, 12, 'sp12_v_b_13')
// (6, 13, 'sp12_v_b_10')
// (6, 14, 'sp12_v_b_9')
// (6, 15, 'sp12_v_b_6')
// (6, 16, 'sp12_v_b_5')
// (6, 17, 'span12_vert_2')
// (7, 6, 'neigh_op_tnl_3')
// (7, 6, 'sp12_h_r_2')
// (7, 7, 'local_g0_3')
// (7, 7, 'local_g1_3')
// (7, 7, 'lutff_2/in_0')
// (7, 7, 'lutff_3/in_2')
// (7, 7, 'neigh_op_lft_3')
// (7, 8, 'neigh_op_bnl_3')
// (8, 6, 'local_g0_5')
// (8, 6, 'local_g1_5')
// (8, 6, 'lutff_0/in_3')
// (8, 6, 'lutff_3/in_3')
// (8, 6, 'sp12_h_r_5')
// (9, 6, 'sp12_h_r_6')
// (10, 6, 'sp12_h_r_9')
// (11, 6, 'sp12_h_r_10')
// (12, 6, 'sp12_h_r_13')
// (13, 6, 'span12_horz_13')

wire n257;
// (5, 6, 'neigh_op_tnr_5')
// (5, 7, 'neigh_op_rgt_5')
// (5, 8, 'neigh_op_bnr_5')
// (6, 6, 'neigh_op_top_5')
// (6, 7, 'local_g1_5')
// (6, 7, 'lutff_2/in_0')
// (6, 7, 'lutff_5/out')
// (6, 7, 'sp4_r_v_b_43')
// (6, 8, 'neigh_op_bot_5')
// (6, 8, 'sp4_r_v_b_30')
// (6, 9, 'sp4_r_v_b_19')
// (6, 10, 'sp4_r_v_b_6')
// (7, 6, 'neigh_op_tnl_5')
// (7, 6, 'sp4_h_r_11')
// (7, 6, 'sp4_v_t_43')
// (7, 7, 'local_g0_5')
// (7, 7, 'local_g1_5')
// (7, 7, 'lutff_2/in_1')
// (7, 7, 'lutff_3/in_3')
// (7, 7, 'neigh_op_lft_5')
// (7, 7, 'sp4_v_b_43')
// (7, 8, 'neigh_op_bnl_5')
// (7, 8, 'sp4_v_b_30')
// (7, 9, 'sp4_v_b_19')
// (7, 10, 'sp4_v_b_6')
// (8, 6, 'local_g0_6')
// (8, 6, 'lutff_1/in_3')
// (8, 6, 'lutff_7/in_3')
// (8, 6, 'sp4_h_r_22')
// (9, 6, 'sp4_h_r_35')
// (10, 6, 'sp4_h_r_46')
// (11, 6, 'sp4_h_l_46')

wire n258;
// (5, 6, 'neigh_op_tnr_6')
// (5, 7, 'neigh_op_rgt_6')
// (5, 8, 'neigh_op_bnr_6')
// (6, 6, 'neigh_op_top_6')
// (6, 7, 'local_g2_6')
// (6, 7, 'lutff_2/in_2')
// (6, 7, 'lutff_6/out')
// (6, 8, 'neigh_op_bot_6')
// (7, 6, 'neigh_op_tnl_6')
// (7, 7, 'local_g0_6')
// (7, 7, 'lutff_5/in_1')
// (7, 7, 'neigh_op_lft_6')
// (7, 8, 'neigh_op_bnl_6')

wire n259;
// (5, 6, 'sp4_r_v_b_39')
// (5, 7, 'sp4_r_v_b_26')
// (5, 8, 'neigh_op_tnr_1')
// (5, 8, 'sp4_r_v_b_15')
// (5, 9, 'neigh_op_rgt_1')
// (5, 9, 'sp4_r_v_b_2')
// (5, 10, 'neigh_op_bnr_1')
// (6, 5, 'sp4_v_t_39')
// (6, 6, 'sp4_v_b_39')
// (6, 7, 'local_g3_2')
// (6, 7, 'lutff_1/in_2')
// (6, 7, 'sp4_v_b_26')
// (6, 8, 'local_g1_1')
// (6, 8, 'lutff_1/in_3')
// (6, 8, 'neigh_op_top_1')
// (6, 8, 'sp4_v_b_15')
// (6, 9, 'lutff_1/out')
// (6, 9, 'sp4_v_b_2')
// (6, 10, 'neigh_op_bot_1')
// (7, 8, 'neigh_op_tnl_1')
// (7, 9, 'neigh_op_lft_1')
// (7, 10, 'neigh_op_bnl_1')

wire n260;
// (5, 7, 'neigh_op_tnr_1')
// (5, 8, 'neigh_op_rgt_1')
// (5, 9, 'neigh_op_bnr_1')
// (6, 6, 'sp4_r_v_b_43')
// (6, 7, 'neigh_op_top_1')
// (6, 7, 'sp4_r_v_b_30')
// (6, 8, 'local_g3_1')
// (6, 8, 'lutff_1/out')
// (6, 8, 'lutff_4/in_0')
// (6, 8, 'sp4_r_v_b_19')
// (6, 9, 'neigh_op_bot_1')
// (6, 9, 'sp4_r_v_b_6')
// (7, 5, 'sp4_v_t_43')
// (7, 6, 'sp4_v_b_43')
// (7, 7, 'local_g3_6')
// (7, 7, 'lutff_4/in_3')
// (7, 7, 'neigh_op_tnl_1')
// (7, 7, 'sp4_v_b_30')
// (7, 8, 'local_g0_1')
// (7, 8, 'local_g0_3')
// (7, 8, 'lutff_2/in_1')
// (7, 8, 'lutff_4/in_3')
// (7, 8, 'lutff_5/in_0')
// (7, 8, 'neigh_op_lft_1')
// (7, 8, 'sp4_v_b_19')
// (7, 9, 'neigh_op_bnl_1')
// (7, 9, 'sp4_v_b_6')

wire n261;
// (5, 7, 'neigh_op_tnr_2')
// (5, 8, 'neigh_op_rgt_2')
// (5, 9, 'neigh_op_bnr_2')
// (6, 7, 'local_g0_2')
// (6, 7, 'local_g1_2')
// (6, 7, 'lutff_3/in_1')
// (6, 7, 'lutff_7/in_2')
// (6, 7, 'neigh_op_top_2')
// (6, 8, 'lutff_2/out')
// (6, 9, 'neigh_op_bot_2')
// (7, 7, 'local_g2_2')
// (7, 7, 'local_g3_2')
// (7, 7, 'lutff_4/in_0')
// (7, 7, 'lutff_6/in_1')
// (7, 7, 'neigh_op_tnl_2')
// (7, 8, 'local_g0_2')
// (7, 8, 'lutff_1/in_1')
// (7, 8, 'lutff_3/in_3')
// (7, 8, 'lutff_5/in_3')
// (7, 8, 'neigh_op_lft_2')
// (7, 9, 'neigh_op_bnl_2')

wire n262;
// (5, 7, 'neigh_op_tnr_3')
// (5, 8, 'neigh_op_rgt_3')
// (5, 9, 'neigh_op_bnr_3')
// (6, 7, 'local_g1_3')
// (6, 7, 'lutff_5/in_1')
// (6, 7, 'neigh_op_top_3')
// (6, 8, 'lutff_3/out')
// (6, 9, 'neigh_op_bot_3')
// (7, 7, 'local_g3_3')
// (7, 7, 'lutff_4/in_2')
// (7, 7, 'neigh_op_tnl_3')
// (7, 8, 'local_g1_3')
// (7, 8, 'lutff_1/in_3')
// (7, 8, 'lutff_3/in_1')
// (7, 8, 'neigh_op_lft_3')
// (7, 9, 'neigh_op_bnl_3')

wire n263;
// (5, 7, 'neigh_op_tnr_4')
// (5, 8, 'neigh_op_rgt_4')
// (5, 9, 'neigh_op_bnr_4')
// (6, 7, 'local_g1_4')
// (6, 7, 'lutff_2/in_3')
// (6, 7, 'neigh_op_top_4')
// (6, 8, 'lutff_4/out')
// (6, 9, 'neigh_op_bot_4')
// (7, 7, 'neigh_op_tnl_4')
// (7, 8, 'neigh_op_lft_4')
// (7, 9, 'neigh_op_bnl_4')

wire n264;
// (5, 7, 'neigh_op_tnr_6')
// (5, 8, 'neigh_op_rgt_6')
// (5, 9, 'neigh_op_bnr_6')
// (6, 7, 'local_g0_6')
// (6, 7, 'local_g1_6')
// (6, 7, 'lutff_1/in_1')
// (6, 7, 'lutff_4/in_3')
// (6, 7, 'lutff_5/in_3')
// (6, 7, 'neigh_op_top_6')
// (6, 8, 'local_g1_6')
// (6, 8, 'lutff_1/in_2')
// (6, 8, 'lutff_6/out')
// (6, 9, 'neigh_op_bot_6')
// (7, 7, 'neigh_op_tnl_6')
// (7, 8, 'neigh_op_lft_6')
// (7, 9, 'neigh_op_bnl_6')

wire n265;
// (5, 7, 'sp4_r_v_b_47')
// (5, 8, 'sp4_r_v_b_34')
// (5, 9, 'sp4_r_v_b_23')
// (5, 10, 'sp4_r_v_b_10')
// (6, 6, 'sp4_v_t_47')
// (6, 7, 'sp4_v_b_47')
// (6, 8, 'sp4_v_b_34')
// (6, 9, 'local_g1_7')
// (6, 9, 'local_g3_0')
// (6, 9, 'lutff_0/in_3')
// (6, 9, 'lutff_1/in_3')
// (6, 9, 'neigh_op_tnr_0')
// (6, 9, 'sp4_v_b_23')
// (6, 10, 'neigh_op_rgt_0')
// (6, 10, 'sp4_h_r_5')
// (6, 10, 'sp4_v_b_10')
// (6, 11, 'neigh_op_bnr_0')
// (7, 9, 'neigh_op_top_0')
// (7, 10, 'lutff_0/out')
// (7, 10, 'sp4_h_r_16')
// (7, 11, 'neigh_op_bot_0')
// (8, 9, 'neigh_op_tnl_0')
// (8, 10, 'neigh_op_lft_0')
// (8, 10, 'sp4_h_r_29')
// (8, 11, 'neigh_op_bnl_0')
// (9, 10, 'sp4_h_r_40')
// (10, 10, 'sp4_h_l_40')

wire n266;
// (5, 8, 'neigh_op_tnr_0')
// (5, 9, 'neigh_op_rgt_0')
// (5, 10, 'neigh_op_bnr_0')
// (6, 6, 'sp4_r_v_b_36')
// (6, 7, 'local_g1_1')
// (6, 7, 'lutff_3/in_3')
// (6, 7, 'sp4_r_v_b_25')
// (6, 8, 'neigh_op_top_0')
// (6, 8, 'sp4_r_v_b_12')
// (6, 9, 'lutff_0/out')
// (6, 9, 'sp4_r_v_b_1')
// (6, 10, 'neigh_op_bot_0')
// (7, 5, 'sp4_v_t_36')
// (7, 6, 'sp4_v_b_36')
// (7, 7, 'local_g2_1')
// (7, 7, 'lutff_6/in_3')
// (7, 7, 'sp4_v_b_25')
// (7, 8, 'neigh_op_tnl_0')
// (7, 8, 'sp4_v_b_12')
// (7, 9, 'neigh_op_lft_0')
// (7, 9, 'sp4_v_b_1')
// (7, 10, 'neigh_op_bnl_0')

wire n267;
// (5, 8, 'neigh_op_tnr_2')
// (5, 9, 'neigh_op_rgt_2')
// (5, 10, 'neigh_op_bnr_2')
// (6, 8, 'neigh_op_top_2')
// (6, 9, 'local_g1_2')
// (6, 9, 'lutff_2/out')
// (6, 9, 'lutff_4/in_3')
// (6, 10, 'neigh_op_bot_2')
// (7, 8, 'neigh_op_tnl_2')
// (7, 9, 'neigh_op_lft_2')
// (7, 10, 'neigh_op_bnl_2')

wire n268;
// (5, 8, 'neigh_op_tnr_3')
// (5, 9, 'neigh_op_rgt_3')
// (5, 10, 'neigh_op_bnr_3')
// (6, 8, 'local_g1_3')
// (6, 8, 'lutff_5/in_3')
// (6, 8, 'neigh_op_top_3')
// (6, 9, 'lutff_3/out')
// (6, 10, 'neigh_op_bot_3')
// (7, 8, 'neigh_op_tnl_3')
// (7, 9, 'neigh_op_lft_3')
// (7, 10, 'neigh_op_bnl_3')

wire n269;
// (5, 8, 'neigh_op_tnr_4')
// (5, 9, 'neigh_op_rgt_4')
// (5, 10, 'neigh_op_bnr_4')
// (6, 8, 'neigh_op_top_4')
// (6, 9, 'local_g0_4')
// (6, 9, 'lutff_3/in_3')
// (6, 9, 'lutff_4/out')
// (6, 10, 'neigh_op_bot_4')
// (7, 8, 'neigh_op_tnl_4')
// (7, 9, 'neigh_op_lft_4')
// (7, 10, 'neigh_op_bnl_4')

wire n270;
// (5, 8, 'neigh_op_tnr_5')
// (5, 9, 'neigh_op_rgt_5')
// (5, 10, 'neigh_op_bnr_5')
// (6, 6, 'sp4_r_v_b_46')
// (6, 7, 'local_g0_0')
// (6, 7, 'local_g2_3')
// (6, 7, 'lutff_4/in_2')
// (6, 7, 'lutff_5/in_2')
// (6, 7, 'sp4_r_v_b_35')
// (6, 8, 'neigh_op_top_5')
// (6, 8, 'sp4_r_v_b_22')
// (6, 9, 'lutff_5/out')
// (6, 9, 'sp4_r_v_b_11')
// (6, 10, 'neigh_op_bot_5')
// (7, 5, 'sp4_v_t_46')
// (7, 6, 'sp4_v_b_46')
// (7, 7, 'sp4_v_b_35')
// (7, 8, 'neigh_op_tnl_5')
// (7, 8, 'sp4_v_b_22')
// (7, 9, 'neigh_op_lft_5')
// (7, 9, 'sp4_v_b_11')
// (7, 10, 'neigh_op_bnl_5')

reg n271 = 0;
// (5, 8, 'neigh_op_tnr_6')
// (5, 9, 'local_g3_6')
// (5, 9, 'lutff_1/in_0')
// (5, 9, 'neigh_op_rgt_6')
// (5, 10, 'neigh_op_bnr_6')
// (6, 8, 'neigh_op_top_6')
// (6, 9, 'lutff_6/out')
// (6, 10, 'neigh_op_bot_6')
// (7, 8, 'neigh_op_tnl_6')
// (7, 9, 'neigh_op_lft_6')
// (7, 10, 'neigh_op_bnl_6')

reg n272 = 0;
// (5, 8, 'neigh_op_tnr_7')
// (5, 9, 'neigh_op_rgt_7')
// (5, 10, 'neigh_op_bnr_7')
// (6, 8, 'neigh_op_top_7')
// (6, 9, 'local_g3_7')
// (6, 9, 'lutff_6/in_0')
// (6, 9, 'lutff_7/out')
// (6, 10, 'neigh_op_bot_7')
// (7, 8, 'neigh_op_tnl_7')
// (7, 9, 'neigh_op_lft_7')
// (7, 10, 'neigh_op_bnl_7')

wire n273;
// (5, 8, 'sp12_h_r_1')
// (6, 8, 'sp12_h_r_2')
// (7, 7, 'neigh_op_tnr_7')
// (7, 8, 'neigh_op_rgt_7')
// (7, 8, 'sp12_h_r_5')
// (7, 9, 'neigh_op_bnr_7')
// (8, 3, 'sp12_v_t_22')
// (8, 4, 'sp12_v_b_22')
// (8, 5, 'sp12_v_b_21')
// (8, 6, 'sp12_v_b_18')
// (8, 7, 'neigh_op_top_7')
// (8, 7, 'sp12_v_b_17')
// (8, 8, 'lutff_7/out')
// (8, 8, 'sp12_h_r_6')
// (8, 8, 'sp12_v_b_14')
// (8, 9, 'neigh_op_bot_7')
// (8, 9, 'sp12_v_b_13')
// (8, 10, 'sp12_v_b_10')
// (8, 11, 'sp12_v_b_9')
// (8, 12, 'local_g2_6')
// (8, 12, 'lutff_0/in_2')
// (8, 12, 'sp12_v_b_6')
// (8, 13, 'sp12_v_b_5')
// (8, 14, 'sp12_v_b_2')
// (8, 15, 'sp12_v_b_1')
// (9, 7, 'neigh_op_tnl_7')
// (9, 8, 'neigh_op_lft_7')
// (9, 8, 'sp12_h_r_9')
// (9, 9, 'neigh_op_bnl_7')
// (10, 8, 'sp12_h_r_10')
// (10, 9, 'sp4_r_v_b_43')
// (10, 10, 'sp4_r_v_b_30')
// (10, 11, 'sp4_r_v_b_19')
// (10, 12, 'sp4_r_v_b_6')
// (11, 8, 'local_g0_5')
// (11, 8, 'lutff_2/in_3')
// (11, 8, 'sp12_h_r_13')
// (11, 8, 'sp4_h_r_6')
// (11, 8, 'sp4_v_t_43')
// (11, 9, 'sp4_v_b_43')
// (11, 10, 'sp4_v_b_30')
// (11, 11, 'sp4_v_b_19')
// (11, 12, 'local_g0_6')
// (11, 12, 'lutff_1/in_3')
// (11, 12, 'lutff_3/in_3')
// (11, 12, 'sp4_v_b_6')
// (12, 8, 'sp12_h_r_14')
// (12, 8, 'sp4_h_r_19')
// (13, 8, 'span12_horz_14')
// (13, 8, 'span4_horz_19')

wire n274;
// (5, 8, 'sp4_h_r_11')
// (6, 8, 'sp4_h_r_22')
// (7, 5, 'neigh_op_tnr_1')
// (7, 6, 'neigh_op_rgt_1')
// (7, 7, 'neigh_op_bnr_1')
// (7, 8, 'sp4_h_r_35')
// (8, 0, 'span12_vert_13')
// (8, 1, 'sp12_v_b_13')
// (8, 2, 'sp12_v_b_10')
// (8, 3, 'sp12_v_b_9')
// (8, 4, 'sp12_v_b_6')
// (8, 5, 'neigh_op_top_1')
// (8, 5, 'sp12_v_b_5')
// (8, 5, 'sp4_r_v_b_46')
// (8, 6, 'lutff_1/out')
// (8, 6, 'sp12_v_b_2')
// (8, 6, 'sp4_r_v_b_35')
// (8, 7, 'local_g3_1')
// (8, 7, 'local_g3_6')
// (8, 7, 'lutff_2/in_0')
// (8, 7, 'lutff_7/in_0')
// (8, 7, 'neigh_op_bot_1')
// (8, 7, 'sp12_v_b_1')
// (8, 7, 'sp4_r_v_b_22')
// (8, 8, 'local_g2_3')
// (8, 8, 'local_g2_6')
// (8, 8, 'lutff_3/in_1')
// (8, 8, 'lutff_7/in_0')
// (8, 8, 'sp4_h_r_46')
// (8, 8, 'sp4_r_v_b_11')
// (9, 4, 'sp4_v_t_46')
// (9, 5, 'neigh_op_tnl_1')
// (9, 5, 'sp4_v_b_46')
// (9, 6, 'neigh_op_lft_1')
// (9, 6, 'sp4_v_b_35')
// (9, 7, 'neigh_op_bnl_1')
// (9, 7, 'sp4_v_b_22')
// (9, 8, 'sp4_h_l_46')
// (9, 8, 'sp4_v_b_11')

wire n275;
// (5, 8, 'sp4_h_r_9')
// (6, 8, 'sp4_h_r_20')
// (7, 7, 'neigh_op_tnr_6')
// (7, 8, 'neigh_op_rgt_6')
// (7, 8, 'sp4_h_r_33')
// (7, 9, 'neigh_op_bnr_6')
// (8, 2, 'sp12_v_t_23')
// (8, 3, 'sp12_v_b_23')
// (8, 4, 'sp12_v_b_20')
// (8, 5, 'sp12_v_b_19')
// (8, 6, 'sp12_v_b_16')
// (8, 7, 'neigh_op_top_6')
// (8, 7, 'sp12_v_b_15')
// (8, 8, 'lutff_6/out')
// (8, 8, 'sp12_v_b_12')
// (8, 8, 'sp4_h_r_44')
// (8, 9, 'neigh_op_bot_6')
// (8, 9, 'sp12_v_b_11')
// (8, 9, 'sp4_r_v_b_39')
// (8, 10, 'sp12_v_b_8')
// (8, 10, 'sp4_r_v_b_26')
// (8, 11, 'sp12_v_b_7')
// (8, 11, 'sp4_r_v_b_15')
// (8, 12, 'sp12_v_b_4')
// (8, 12, 'sp4_r_v_b_2')
// (8, 13, 'local_g3_3')
// (8, 13, 'lutff_3/in_3')
// (8, 13, 'lutff_4/in_2')
// (8, 13, 'sp12_v_b_3')
// (8, 14, 'sp12_v_b_0')
// (9, 7, 'neigh_op_tnl_6')
// (9, 8, 'local_g1_6')
// (9, 8, 'lutff_5/in_2')
// (9, 8, 'neigh_op_lft_6')
// (9, 8, 'sp4_h_l_44')
// (9, 8, 'sp4_v_t_39')
// (9, 9, 'neigh_op_bnl_6')
// (9, 9, 'sp4_v_b_39')
// (9, 10, 'sp4_v_b_26')
// (9, 11, 'sp4_v_b_15')
// (9, 12, 'local_g0_2')
// (9, 12, 'lutff_7/in_3')
// (9, 12, 'sp4_h_r_8')
// (9, 12, 'sp4_v_b_2')
// (10, 12, 'sp4_h_r_21')
// (11, 12, 'local_g3_0')
// (11, 12, 'lutff_6/in_3')
// (11, 12, 'lutff_7/in_2')
// (11, 12, 'sp4_h_r_32')
// (12, 12, 'sp4_h_r_45')
// (13, 12, 'span4_horz_45')

wire n276;
// (5, 8, 'sp4_r_v_b_36')
// (5, 9, 'sp4_r_v_b_25')
// (5, 10, 'sp4_r_v_b_12')
// (5, 11, 'neigh_op_tnr_4')
// (5, 11, 'sp4_r_v_b_1')
// (5, 12, 'neigh_op_rgt_4')
// (5, 12, 'sp4_r_v_b_40')
// (5, 13, 'neigh_op_bnr_4')
// (5, 13, 'sp4_r_v_b_29')
// (5, 14, 'sp4_r_v_b_16')
// (5, 15, 'sp4_r_v_b_5')
// (6, 4, 'sp12_v_t_23')
// (6, 5, 'sp12_v_b_23')
// (6, 5, 'sp4_r_v_b_40')
// (6, 6, 'sp12_v_b_20')
// (6, 6, 'sp4_r_v_b_29')
// (6, 7, 'local_g3_3')
// (6, 7, 'lutff_1/in_3')
// (6, 7, 'sp12_v_b_19')
// (6, 7, 'sp4_h_r_1')
// (6, 7, 'sp4_r_v_b_16')
// (6, 7, 'sp4_v_t_36')
// (6, 8, 'local_g2_0')
// (6, 8, 'local_g3_0')
// (6, 8, 'lutff_2/in_2')
// (6, 8, 'lutff_3/in_2')
// (6, 8, 'lutff_5/in_2')
// (6, 8, 'lutff_6/in_2')
// (6, 8, 'lutff_7/in_3')
// (6, 8, 'sp12_v_b_16')
// (6, 8, 'sp4_r_v_b_5')
// (6, 8, 'sp4_v_b_36')
// (6, 9, 'local_g2_7')
// (6, 9, 'lutff_0/in_1')
// (6, 9, 'sp12_v_b_15')
// (6, 9, 'sp4_r_v_b_44')
// (6, 9, 'sp4_v_b_25')
// (6, 10, 'sp12_v_b_12')
// (6, 10, 'sp4_r_v_b_33')
// (6, 10, 'sp4_v_b_12')
// (6, 11, 'neigh_op_top_4')
// (6, 11, 'sp12_v_b_11')
// (6, 11, 'sp4_r_v_b_20')
// (6, 11, 'sp4_v_b_1')
// (6, 11, 'sp4_v_t_40')
// (6, 12, 'lutff_4/out')
// (6, 12, 'sp12_v_b_8')
// (6, 12, 'sp4_r_v_b_9')
// (6, 12, 'sp4_v_b_40')
// (6, 13, 'neigh_op_bot_4')
// (6, 13, 'sp12_v_b_7')
// (6, 13, 'sp4_v_b_29')
// (6, 14, 'sp12_v_b_4')
// (6, 14, 'sp4_v_b_16')
// (6, 15, 'sp12_v_b_3')
// (6, 15, 'sp4_v_b_5')
// (6, 16, 'sp12_v_b_0')
// (7, 4, 'sp4_v_t_40')
// (7, 5, 'sp4_v_b_40')
// (7, 6, 'sp4_v_b_29')
// (7, 7, 'local_g0_0')
// (7, 7, 'lutff_0/in_2')
// (7, 7, 'sp4_h_r_12')
// (7, 7, 'sp4_v_b_16')
// (7, 8, 'local_g0_5')
// (7, 8, 'lutff_5/in_2')
// (7, 8, 'sp4_v_b_5')
// (7, 8, 'sp4_v_t_44')
// (7, 9, 'sp4_v_b_44')
// (7, 10, 'sp4_v_b_33')
// (7, 11, 'neigh_op_tnl_4')
// (7, 11, 'sp4_v_b_20')
// (7, 12, 'neigh_op_lft_4')
// (7, 12, 'sp4_v_b_9')
// (7, 13, 'neigh_op_bnl_4')
// (8, 7, 'local_g2_1')
// (8, 7, 'lutff_4/in_3')
// (8, 7, 'lutff_6/in_1')
// (8, 7, 'sp4_h_r_25')
// (9, 7, 'sp4_h_r_36')
// (10, 7, 'sp4_h_l_36')

reg n277 = 0;
// (5, 9, 'neigh_op_tnr_0')
// (5, 10, 'neigh_op_rgt_0')
// (5, 11, 'neigh_op_bnr_0')
// (6, 9, 'neigh_op_top_0')
// (6, 10, 'lutff_0/out')
// (6, 11, 'neigh_op_bot_0')
// (7, 9, 'neigh_op_tnl_0')
// (7, 10, 'local_g0_0')
// (7, 10, 'lutff_3/in_1')
// (7, 10, 'lutff_7/in_1')
// (7, 10, 'neigh_op_lft_0')
// (7, 11, 'neigh_op_bnl_0')

reg n278 = 0;
// (5, 9, 'neigh_op_tnr_1')
// (5, 10, 'neigh_op_rgt_1')
// (5, 11, 'neigh_op_bnr_1')
// (6, 9, 'neigh_op_top_1')
// (6, 10, 'local_g1_1')
// (6, 10, 'lutff_1/out')
// (6, 10, 'lutff_6/in_0')
// (6, 11, 'neigh_op_bot_1')
// (7, 9, 'neigh_op_tnl_1')
// (7, 10, 'neigh_op_lft_1')
// (7, 11, 'neigh_op_bnl_1')

reg n279 = 0;
// (5, 9, 'neigh_op_tnr_2')
// (5, 10, 'neigh_op_rgt_2')
// (5, 11, 'neigh_op_bnr_2')
// (6, 9, 'neigh_op_top_2')
// (6, 10, 'lutff_2/out')
// (6, 11, 'neigh_op_bot_2')
// (7, 9, 'neigh_op_tnl_2')
// (7, 10, 'local_g0_2')
// (7, 10, 'lutff_6/in_0')
// (7, 10, 'neigh_op_lft_2')
// (7, 11, 'neigh_op_bnl_2')

reg n280 = 0;
// (5, 9, 'neigh_op_tnr_3')
// (5, 10, 'neigh_op_rgt_3')
// (5, 11, 'neigh_op_bnr_3')
// (6, 9, 'neigh_op_top_3')
// (6, 10, 'local_g0_3')
// (6, 10, 'lutff_3/out')
// (6, 10, 'lutff_5/in_0')
// (6, 11, 'neigh_op_bot_3')
// (7, 9, 'neigh_op_tnl_3')
// (7, 10, 'neigh_op_lft_3')
// (7, 11, 'neigh_op_bnl_3')

reg n281 = 0;
// (5, 9, 'neigh_op_tnr_4')
// (5, 10, 'neigh_op_rgt_4')
// (5, 11, 'neigh_op_bnr_4')
// (6, 9, 'neigh_op_top_4')
// (6, 10, 'local_g1_4')
// (6, 10, 'lutff_3/in_0')
// (6, 10, 'lutff_4/out')
// (6, 11, 'neigh_op_bot_4')
// (7, 9, 'neigh_op_tnl_4')
// (7, 10, 'neigh_op_lft_4')
// (7, 11, 'neigh_op_bnl_4')

reg n282 = 0;
// (5, 9, 'neigh_op_tnr_5')
// (5, 10, 'neigh_op_rgt_5')
// (5, 11, 'neigh_op_bnr_5')
// (6, 9, 'neigh_op_top_5')
// (6, 10, 'local_g1_5')
// (6, 10, 'lutff_2/in_0')
// (6, 10, 'lutff_5/out')
// (6, 11, 'neigh_op_bot_5')
// (7, 9, 'neigh_op_tnl_5')
// (7, 10, 'neigh_op_lft_5')
// (7, 11, 'neigh_op_bnl_5')

reg n283 = 0;
// (5, 9, 'neigh_op_tnr_6')
// (5, 10, 'neigh_op_rgt_6')
// (5, 11, 'neigh_op_bnr_6')
// (6, 9, 'neigh_op_top_6')
// (6, 10, 'local_g0_6')
// (6, 10, 'lutff_0/in_0')
// (6, 10, 'lutff_6/out')
// (6, 11, 'neigh_op_bot_6')
// (7, 9, 'neigh_op_tnl_6')
// (7, 10, 'neigh_op_lft_6')
// (7, 11, 'neigh_op_bnl_6')

reg n284 = 0;
// (5, 9, 'neigh_op_tnr_7')
// (5, 10, 'neigh_op_rgt_7')
// (5, 11, 'neigh_op_bnr_7')
// (6, 9, 'neigh_op_top_7')
// (6, 10, 'local_g1_7')
// (6, 10, 'lutff_4/in_0')
// (6, 10, 'lutff_7/out')
// (6, 11, 'neigh_op_bot_7')
// (7, 9, 'neigh_op_tnl_7')
// (7, 10, 'neigh_op_lft_7')
// (7, 11, 'neigh_op_bnl_7')

wire n285;
// (5, 9, 'sp4_r_v_b_37')
// (5, 10, 'sp4_r_v_b_24')
// (5, 11, 'neigh_op_tnr_0')
// (5, 11, 'sp4_r_v_b_13')
// (5, 12, 'neigh_op_rgt_0')
// (5, 12, 'sp4_r_v_b_0')
// (5, 13, 'neigh_op_bnr_0')
// (6, 8, 'sp4_v_t_37')
// (6, 9, 'sp4_v_b_37')
// (6, 10, 'sp4_v_b_24')
// (6, 11, 'local_g1_5')
// (6, 11, 'lutff_1/in_3')
// (6, 11, 'neigh_op_top_0')
// (6, 11, 'sp4_v_b_13')
// (6, 12, 'lutff_0/out')
// (6, 12, 'sp4_v_b_0')
// (6, 13, 'neigh_op_bot_0')
// (7, 11, 'neigh_op_tnl_0')
// (7, 12, 'neigh_op_lft_0')
// (7, 13, 'neigh_op_bnl_0')

wire n286;
// (5, 10, 'local_g2_2')
// (5, 10, 'lutff_2/in_0')
// (5, 10, 'lutff_7/in_3')
// (5, 10, 'neigh_op_tnr_2')
// (5, 11, 'neigh_op_rgt_2')
// (5, 12, 'local_g1_2')
// (5, 12, 'lutff_2/in_3')
// (5, 12, 'neigh_op_bnr_2')
// (6, 8, 'sp4_r_v_b_40')
// (6, 9, 'local_g0_5')
// (6, 9, 'local_g1_5')
// (6, 9, 'lutff_3/in_0')
// (6, 9, 'lutff_7/in_3')
// (6, 9, 'sp4_r_v_b_29')
// (6, 10, 'neigh_op_top_2')
// (6, 10, 'sp4_r_v_b_16')
// (6, 11, 'local_g1_2')
// (6, 11, 'local_g2_2')
// (6, 11, 'lutff_0/in_0')
// (6, 11, 'lutff_1/in_0')
// (6, 11, 'lutff_2/out')
// (6, 11, 'lutff_4/in_3')
// (6, 11, 'sp4_r_v_b_37')
// (6, 11, 'sp4_r_v_b_5')
// (6, 12, 'local_g0_2')
// (6, 12, 'lutff_4/in_0')
// (6, 12, 'lutff_5/in_3')
// (6, 12, 'neigh_op_bot_2')
// (6, 12, 'sp4_r_v_b_24')
// (6, 13, 'sp4_r_v_b_13')
// (6, 14, 'sp4_r_v_b_0')
// (7, 7, 'sp4_v_t_40')
// (7, 8, 'sp4_v_b_40')
// (7, 9, 'sp4_v_b_29')
// (7, 10, 'local_g2_2')
// (7, 10, 'lutff_0/in_0')
// (7, 10, 'lutff_4/in_0')
// (7, 10, 'lutff_5/in_3')
// (7, 10, 'neigh_op_tnl_2')
// (7, 10, 'sp4_v_b_16')
// (7, 10, 'sp4_v_t_37')
// (7, 11, 'local_g1_2')
// (7, 11, 'lutff_1/in_0')
// (7, 11, 'neigh_op_lft_2')
// (7, 11, 'sp4_v_b_37')
// (7, 11, 'sp4_v_b_5')
// (7, 12, 'local_g2_2')
// (7, 12, 'lutff_5/in_3')
// (7, 12, 'neigh_op_bnl_2')
// (7, 12, 'sp4_v_b_24')
// (7, 13, 'local_g0_5')
// (7, 13, 'lutff_0/in_3')
// (7, 13, 'sp4_v_b_13')
// (7, 14, 'sp4_v_b_0')

wire n287;
// (5, 10, 'neigh_op_tnr_0')
// (5, 11, 'neigh_op_rgt_0')
// (5, 12, 'neigh_op_bnr_0')
// (6, 0, 'span12_vert_20')
// (6, 1, 'sp12_v_b_20')
// (6, 2, 'sp12_v_b_19')
// (6, 3, 'sp12_v_b_16')
// (6, 4, 'sp12_v_b_15')
// (6, 5, 'sp12_v_b_12')
// (6, 6, 'sp12_v_b_11')
// (6, 7, 'sp12_v_b_8')
// (6, 8, 'local_g2_7')
// (6, 8, 'local_g3_7')
// (6, 8, 'lutff_2/in_1')
// (6, 8, 'lutff_3/in_1')
// (6, 8, 'lutff_5/in_1')
// (6, 8, 'lutff_6/in_1')
// (6, 8, 'lutff_7/in_2')
// (6, 8, 'sp12_v_b_7')
// (6, 9, 'sp12_v_b_4')
// (6, 10, 'neigh_op_top_0')
// (6, 10, 'sp12_v_b_3')
// (6, 11, 'lutff_0/out')
// (6, 11, 'sp12_v_b_0')
// (6, 12, 'neigh_op_bot_0')
// (7, 10, 'neigh_op_tnl_0')
// (7, 11, 'neigh_op_lft_0')
// (7, 12, 'neigh_op_bnl_0')

wire n288;
// (5, 10, 'neigh_op_tnr_1')
// (5, 11, 'neigh_op_rgt_1')
// (5, 12, 'neigh_op_bnr_1')
// (6, 0, 'span12_vert_22')
// (6, 1, 'sp12_v_b_22')
// (6, 2, 'sp12_v_b_21')
// (6, 3, 'sp12_v_b_18')
// (6, 4, 'sp12_v_b_17')
// (6, 5, 'sp12_v_b_14')
// (6, 6, 'sp12_v_b_13')
// (6, 7, 'sp12_v_b_10')
// (6, 8, 'local_g2_1')
// (6, 8, 'lutff_2/in_3')
// (6, 8, 'lutff_4/in_1')
// (6, 8, 'sp12_v_b_9')
// (6, 9, 'local_g3_6')
// (6, 9, 'lutff_5/in_2')
// (6, 9, 'sp12_v_b_6')
// (6, 10, 'neigh_op_top_1')
// (6, 10, 'sp12_v_b_5')
// (6, 11, 'lutff_1/out')
// (6, 11, 'sp12_v_b_2')
// (6, 12, 'neigh_op_bot_1')
// (6, 12, 'sp12_v_b_1')
// (7, 10, 'neigh_op_tnl_1')
// (7, 11, 'neigh_op_lft_1')
// (7, 12, 'neigh_op_bnl_1')

reg n289 = 0;
// (5, 10, 'neigh_op_tnr_3')
// (5, 11, 'neigh_op_rgt_3')
// (5, 12, 'neigh_op_bnr_3')
// (6, 10, 'neigh_op_top_3')
// (6, 11, 'lutff_3/out')
// (6, 12, 'local_g0_3')
// (6, 12, 'lutff_7/in_0')
// (6, 12, 'neigh_op_bot_3')
// (7, 10, 'neigh_op_tnl_3')
// (7, 11, 'neigh_op_lft_3')
// (7, 12, 'neigh_op_bnl_3')

reg n290 = 0;
// (5, 10, 'neigh_op_tnr_4')
// (5, 11, 'neigh_op_rgt_4')
// (5, 12, 'neigh_op_bnr_4')
// (6, 10, 'neigh_op_top_4')
// (6, 11, 'local_g1_4')
// (6, 11, 'lutff_4/out')
// (6, 11, 'lutff_7/in_0')
// (6, 12, 'neigh_op_bot_4')
// (7, 10, 'neigh_op_tnl_4')
// (7, 11, 'neigh_op_lft_4')
// (7, 12, 'neigh_op_bnl_4')

reg n291 = 0;
// (5, 10, 'neigh_op_tnr_7')
// (5, 11, 'neigh_op_rgt_7')
// (5, 12, 'neigh_op_bnr_7')
// (6, 10, 'neigh_op_top_7')
// (6, 11, 'local_g0_7')
// (6, 11, 'lutff_3/in_0')
// (6, 11, 'lutff_7/out')
// (6, 12, 'neigh_op_bot_7')
// (7, 10, 'neigh_op_tnl_7')
// (7, 11, 'neigh_op_lft_7')
// (7, 12, 'neigh_op_bnl_7')

wire n292;
// (5, 11, 'neigh_op_tnr_2')
// (5, 12, 'neigh_op_rgt_2')
// (5, 13, 'neigh_op_bnr_2')
// (6, 11, 'neigh_op_top_2')
// (6, 12, 'local_g2_2')
// (6, 12, 'lutff_2/out')
// (6, 12, 'lutff_3/in_3')
// (6, 13, 'neigh_op_bot_2')
// (7, 11, 'neigh_op_tnl_2')
// (7, 12, 'neigh_op_lft_2')
// (7, 13, 'neigh_op_bnl_2')

wire n293;
// (5, 11, 'neigh_op_tnr_3')
// (5, 12, 'neigh_op_rgt_3')
// (5, 13, 'neigh_op_bnr_3')
// (6, 3, 'sp12_v_t_22')
// (6, 4, 'sp12_v_b_22')
// (6, 5, 'sp12_v_b_21')
// (6, 6, 'sp12_v_b_18')
// (6, 7, 'sp12_v_b_17')
// (6, 8, 'sp12_v_b_14')
// (6, 9, 'sp12_v_b_13')
// (6, 10, 'sp12_v_b_10')
// (6, 11, 'local_g2_1')
// (6, 11, 'lutff_0/in_3')
// (6, 11, 'neigh_op_top_3')
// (6, 11, 'sp12_v_b_9')
// (6, 12, 'lutff_3/out')
// (6, 12, 'sp12_v_b_6')
// (6, 13, 'neigh_op_bot_3')
// (6, 13, 'sp12_v_b_5')
// (6, 14, 'sp12_v_b_2')
// (6, 15, 'sp12_v_b_1')
// (7, 11, 'neigh_op_tnl_3')
// (7, 12, 'neigh_op_lft_3')
// (7, 13, 'neigh_op_bnl_3')

reg n294 = 0;
// (5, 11, 'neigh_op_tnr_5')
// (5, 12, 'local_g2_5')
// (5, 12, 'lutff_7/in_0')
// (5, 12, 'neigh_op_rgt_5')
// (5, 13, 'neigh_op_bnr_5')
// (6, 11, 'neigh_op_top_5')
// (6, 12, 'lutff_5/out')
// (6, 13, 'neigh_op_bot_5')
// (7, 11, 'neigh_op_tnl_5')
// (7, 12, 'neigh_op_lft_5')
// (7, 13, 'neigh_op_bnl_5')

reg n295 = 0;
// (5, 11, 'neigh_op_tnr_7')
// (5, 12, 'neigh_op_rgt_7')
// (5, 13, 'neigh_op_bnr_7')
// (6, 11, 'neigh_op_top_7')
// (6, 12, 'local_g0_7')
// (6, 12, 'lutff_2/in_1')
// (6, 12, 'lutff_6/in_1')
// (6, 12, 'lutff_7/out')
// (6, 13, 'neigh_op_bot_7')
// (7, 11, 'neigh_op_tnl_7')
// (7, 12, 'neigh_op_lft_7')
// (7, 13, 'neigh_op_bnl_7')

reg n296 = 0;
// (5, 12, 'neigh_op_tnr_0')
// (5, 13, 'neigh_op_rgt_0')
// (5, 14, 'neigh_op_bnr_0')
// (6, 11, 'sp4_r_v_b_41')
// (6, 12, 'local_g0_4')
// (6, 12, 'local_g1_4')
// (6, 12, 'lutff_0/in_0')
// (6, 12, 'lutff_5/in_0')
// (6, 12, 'neigh_op_top_0')
// (6, 12, 'sp4_r_v_b_28')
// (6, 13, 'local_g0_0')
// (6, 13, 'local_g1_0')
// (6, 13, 'lutff_0/out')
// (6, 13, 'lutff_6/in_0')
// (6, 13, 'lutff_7/in_0')
// (6, 13, 'sp4_r_v_b_17')
// (6, 14, 'neigh_op_bot_0')
// (6, 14, 'sp4_r_v_b_4')
// (7, 10, 'sp4_v_t_41')
// (7, 11, 'sp4_v_b_41')
// (7, 12, 'neigh_op_tnl_0')
// (7, 12, 'sp4_v_b_28')
// (7, 13, 'neigh_op_lft_0')
// (7, 13, 'sp4_v_b_17')
// (7, 14, 'neigh_op_bnl_0')
// (7, 14, 'sp4_v_b_4')

reg n297 = 0;
// (5, 12, 'neigh_op_tnr_1')
// (5, 13, 'neigh_op_rgt_1')
// (5, 14, 'neigh_op_bnr_1')
// (6, 12, 'neigh_op_top_1')
// (6, 13, 'local_g1_1')
// (6, 13, 'lutff_1/out')
// (6, 13, 'lutff_2/in_0')
// (6, 14, 'neigh_op_bot_1')
// (7, 12, 'neigh_op_tnl_1')
// (7, 13, 'neigh_op_lft_1')
// (7, 14, 'neigh_op_bnl_1')

reg n298 = 0;
// (5, 12, 'neigh_op_tnr_2')
// (5, 13, 'local_g1_1')
// (5, 13, 'lutff_0/in_0')
// (5, 13, 'neigh_op_rgt_2')
// (5, 13, 'sp4_h_r_9')
// (5, 14, 'neigh_op_bnr_2')
// (6, 12, 'neigh_op_top_2')
// (6, 13, 'local_g0_2')
// (6, 13, 'lutff_2/out')
// (6, 13, 'lutff_7/in_1')
// (6, 13, 'sp4_h_r_20')
// (6, 14, 'neigh_op_bot_2')
// (7, 12, 'neigh_op_tnl_2')
// (7, 13, 'neigh_op_lft_2')
// (7, 13, 'sp4_h_r_33')
// (7, 14, 'neigh_op_bnl_2')
// (8, 13, 'sp4_h_r_44')
// (9, 13, 'sp4_h_l_44')

reg n299 = 0;
// (5, 12, 'neigh_op_tnr_3')
// (5, 13, 'neigh_op_rgt_3')
// (5, 14, 'neigh_op_bnr_3')
// (6, 12, 'neigh_op_top_3')
// (6, 13, 'local_g1_3')
// (6, 13, 'lutff_0/in_0')
// (6, 13, 'lutff_3/out')
// (6, 14, 'neigh_op_bot_3')
// (7, 12, 'neigh_op_tnl_3')
// (7, 13, 'neigh_op_lft_3')
// (7, 14, 'neigh_op_bnl_3')

reg n300 = 0;
// (5, 12, 'neigh_op_tnr_4')
// (5, 13, 'neigh_op_rgt_4')
// (5, 14, 'neigh_op_bnr_4')
// (6, 12, 'neigh_op_top_4')
// (6, 13, 'local_g1_4')
// (6, 13, 'lutff_1/in_0')
// (6, 13, 'lutff_4/out')
// (6, 14, 'neigh_op_bot_4')
// (7, 12, 'neigh_op_tnl_4')
// (7, 13, 'neigh_op_lft_4')
// (7, 14, 'neigh_op_bnl_4')

reg n301 = 0;
// (5, 12, 'neigh_op_tnr_5')
// (5, 13, 'neigh_op_rgt_5')
// (5, 14, 'neigh_op_bnr_5')
// (6, 12, 'neigh_op_top_5')
// (6, 13, 'local_g0_5')
// (6, 13, 'lutff_3/in_0')
// (6, 13, 'lutff_5/out')
// (6, 14, 'neigh_op_bot_5')
// (7, 12, 'neigh_op_tnl_5')
// (7, 13, 'neigh_op_lft_5')
// (7, 14, 'neigh_op_bnl_5')

reg n302 = 0;
// (5, 12, 'neigh_op_tnr_6')
// (5, 13, 'neigh_op_rgt_6')
// (5, 14, 'neigh_op_bnr_6')
// (6, 12, 'neigh_op_top_6')
// (6, 13, 'local_g0_6')
// (6, 13, 'lutff_4/in_0')
// (6, 13, 'lutff_6/out')
// (6, 14, 'neigh_op_bot_6')
// (7, 12, 'neigh_op_tnl_6')
// (7, 13, 'neigh_op_lft_6')
// (7, 14, 'neigh_op_bnl_6')

reg n303 = 0;
// (5, 12, 'neigh_op_tnr_7')
// (5, 13, 'neigh_op_rgt_7')
// (5, 14, 'neigh_op_bnr_7')
// (6, 12, 'neigh_op_top_7')
// (6, 13, 'local_g0_7')
// (6, 13, 'lutff_5/in_0')
// (6, 13, 'lutff_7/out')
// (6, 14, 'neigh_op_bot_7')
// (7, 12, 'neigh_op_tnl_7')
// (7, 13, 'neigh_op_lft_7')
// (7, 14, 'neigh_op_bnl_7')

wire n304;
// (6, 1, 'neigh_op_tnr_0')
// (6, 2, 'neigh_op_rgt_0')
// (6, 3, 'neigh_op_bnr_0')
// (7, 1, 'neigh_op_top_0')
// (7, 2, 'local_g2_0')
// (7, 2, 'local_g3_0')
// (7, 2, 'lutff_0/out')
// (7, 2, 'lutff_4/in_2')
// (7, 2, 'lutff_7/in_2')
// (7, 3, 'neigh_op_bot_0')
// (8, 1, 'neigh_op_tnl_0')
// (8, 2, 'neigh_op_lft_0')
// (8, 3, 'neigh_op_bnl_0')

wire n305;
// (6, 1, 'neigh_op_tnr_1')
// (6, 2, 'neigh_op_rgt_1')
// (6, 3, 'neigh_op_bnr_1')
// (7, 1, 'neigh_op_top_1')
// (7, 2, 'lutff_1/out')
// (7, 3, 'neigh_op_bot_1')
// (8, 1, 'neigh_op_tnl_1')
// (8, 2, 'neigh_op_lft_1')
// (8, 3, 'local_g2_1')
// (8, 3, 'lutff_4/in_3')
// (8, 3, 'lutff_6/in_3')
// (8, 3, 'neigh_op_bnl_1')

wire n306;
// (6, 1, 'neigh_op_tnr_2')
// (6, 2, 'neigh_op_rgt_2')
// (6, 3, 'neigh_op_bnr_2')
// (7, 1, 'neigh_op_top_2')
// (7, 2, 'local_g2_2')
// (7, 2, 'lutff_1/in_1')
// (7, 2, 'lutff_2/out')
// (7, 2, 'lutff_3/in_1')
// (7, 3, 'neigh_op_bot_2')
// (8, 1, 'neigh_op_tnl_2')
// (8, 2, 'local_g0_2')
// (8, 2, 'local_g1_2')
// (8, 2, 'lutff_1/in_1')
// (8, 2, 'lutff_2/in_3')
// (8, 2, 'lutff_3/in_0')
// (8, 2, 'lutff_4/in_1')
// (8, 2, 'lutff_5/in_2')
// (8, 2, 'lutff_6/in_2')
// (8, 2, 'lutff_7/in_0')
// (8, 2, 'neigh_op_lft_2')
// (8, 3, 'neigh_op_bnl_2')

wire n307;
// (6, 1, 'neigh_op_tnr_3')
// (6, 2, 'neigh_op_rgt_3')
// (6, 2, 'sp4_r_v_b_38')
// (6, 3, 'neigh_op_bnr_3')
// (6, 3, 'sp4_r_v_b_27')
// (6, 4, 'sp4_r_v_b_14')
// (6, 5, 'sp4_r_v_b_3')
// (7, 1, 'neigh_op_top_3')
// (7, 1, 'sp4_v_t_38')
// (7, 2, 'lutff_3/out')
// (7, 2, 'sp4_r_v_b_39')
// (7, 2, 'sp4_v_b_38')
// (7, 3, 'neigh_op_bot_3')
// (7, 3, 'sp4_r_v_b_26')
// (7, 3, 'sp4_v_b_27')
// (7, 4, 'local_g0_6')
// (7, 4, 'lutff_1/in_3')
// (7, 4, 'sp4_r_v_b_15')
// (7, 4, 'sp4_v_b_14')
// (7, 5, 'sp4_r_v_b_2')
// (7, 5, 'sp4_v_b_3')
// (8, 1, 'neigh_op_tnl_3')
// (8, 1, 'sp4_v_t_39')
// (8, 2, 'neigh_op_lft_3')
// (8, 2, 'sp4_v_b_39')
// (8, 3, 'neigh_op_bnl_3')
// (8, 3, 'sp4_v_b_26')
// (8, 4, 'local_g0_7')
// (8, 4, 'lutff_2/in_3')
// (8, 4, 'sp4_v_b_15')
// (8, 5, 'sp4_v_b_2')

wire n308;
// (6, 1, 'neigh_op_tnr_4')
// (6, 2, 'neigh_op_rgt_4')
// (6, 3, 'neigh_op_bnr_4')
// (7, 1, 'neigh_op_top_4')
// (7, 2, 'lutff_4/out')
// (7, 3, 'neigh_op_bot_4')
// (8, 1, 'neigh_op_tnl_4')
// (8, 2, 'local_g0_4')
// (8, 2, 'local_g1_4')
// (8, 2, 'lutff_1/in_0')
// (8, 2, 'lutff_2/in_2')
// (8, 2, 'lutff_3/in_2')
// (8, 2, 'lutff_4/in_3')
// (8, 2, 'lutff_5/in_0')
// (8, 2, 'lutff_6/in_0')
// (8, 2, 'lutff_7/in_1')
// (8, 2, 'neigh_op_lft_4')
// (8, 3, 'neigh_op_bnl_4')

wire n309;
// (6, 1, 'neigh_op_tnr_5')
// (6, 2, 'neigh_op_rgt_5')
// (6, 3, 'neigh_op_bnr_5')
// (7, 1, 'neigh_op_top_5')
// (7, 2, 'local_g0_5')
// (7, 2, 'lutff_1/in_2')
// (7, 2, 'lutff_3/in_2')
// (7, 2, 'lutff_5/out')
// (7, 3, 'neigh_op_bot_5')
// (8, 1, 'neigh_op_tnl_5')
// (8, 2, 'neigh_op_lft_5')
// (8, 3, 'neigh_op_bnl_5')

wire n310;
// (6, 1, 'neigh_op_tnr_6')
// (6, 2, 'neigh_op_rgt_6')
// (6, 3, 'neigh_op_bnr_6')
// (7, 1, 'neigh_op_top_6')
// (7, 2, 'local_g1_6')
// (7, 2, 'lutff_5/in_2')
// (7, 2, 'lutff_6/out')
// (7, 3, 'neigh_op_bot_6')
// (8, 1, 'neigh_op_tnl_6')
// (8, 2, 'local_g1_6')
// (8, 2, 'lutff_0/in_3')
// (8, 2, 'neigh_op_lft_6')
// (8, 3, 'neigh_op_bnl_6')

wire n311;
// (6, 1, 'neigh_op_tnr_7')
// (6, 2, 'neigh_op_rgt_7')
// (6, 3, 'neigh_op_bnr_7')
// (7, 1, 'neigh_op_top_7')
// (7, 2, 'local_g0_7')
// (7, 2, 'lutff_1/in_0')
// (7, 2, 'lutff_3/in_0')
// (7, 2, 'lutff_7/out')
// (7, 3, 'neigh_op_bot_7')
// (8, 1, 'neigh_op_tnl_7')
// (8, 2, 'local_g0_7')
// (8, 2, 'lutff_7/in_2')
// (8, 2, 'neigh_op_lft_7')
// (8, 3, 'neigh_op_bnl_7')

wire n312;
// (6, 1, 'sp4_r_v_b_36')
// (6, 2, 'neigh_op_tnr_6')
// (6, 2, 'sp4_r_v_b_25')
// (6, 3, 'neigh_op_rgt_6')
// (6, 3, 'sp4_r_v_b_12')
// (6, 4, 'neigh_op_bnr_6')
// (6, 4, 'sp4_r_v_b_1')
// (7, 0, 'span4_vert_36')
// (7, 1, 'sp4_v_b_36')
// (7, 2, 'local_g2_1')
// (7, 2, 'lutff_5/in_0')
// (7, 2, 'lutff_7/in_0')
// (7, 2, 'neigh_op_top_6')
// (7, 2, 'sp4_v_b_25')
// (7, 3, 'lutff_6/out')
// (7, 3, 'sp4_v_b_12')
// (7, 4, 'neigh_op_bot_6')
// (7, 4, 'sp4_v_b_1')
// (8, 2, 'local_g2_6')
// (8, 2, 'local_g3_6')
// (8, 2, 'lutff_1/in_2')
// (8, 2, 'lutff_2/in_0')
// (8, 2, 'lutff_3/in_3')
// (8, 2, 'lutff_4/in_2')
// (8, 2, 'lutff_5/in_1')
// (8, 2, 'lutff_6/in_1')
// (8, 2, 'neigh_op_tnl_6')
// (8, 3, 'neigh_op_lft_6')
// (8, 4, 'neigh_op_bnl_6')

wire n313;
// (6, 1, 'sp4_r_v_b_38')
// (6, 2, 'neigh_op_tnr_7')
// (6, 2, 'sp4_r_v_b_27')
// (6, 3, 'neigh_op_rgt_7')
// (6, 3, 'sp4_r_v_b_14')
// (6, 4, 'neigh_op_bnr_7')
// (6, 4, 'sp4_r_v_b_3')
// (7, 0, 'span4_vert_38')
// (7, 1, 'sp4_v_b_38')
// (7, 2, 'local_g2_3')
// (7, 2, 'lutff_6/in_3')
// (7, 2, 'neigh_op_top_7')
// (7, 2, 'sp4_v_b_27')
// (7, 3, 'lutff_7/out')
// (7, 3, 'sp4_v_b_14')
// (7, 4, 'neigh_op_bot_7')
// (7, 4, 'sp4_v_b_3')
// (8, 2, 'neigh_op_tnl_7')
// (8, 3, 'neigh_op_lft_7')
// (8, 4, 'neigh_op_bnl_7')

wire n314;
// (6, 1, 'sp4_r_v_b_40')
// (6, 2, 'sp4_r_v_b_29')
// (6, 3, 'local_g3_3')
// (6, 3, 'lutff_6/in_2')
// (6, 3, 'neigh_op_tnr_3')
// (6, 3, 'sp4_r_v_b_16')
// (6, 4, 'neigh_op_rgt_3')
// (6, 4, 'sp4_r_v_b_5')
// (6, 5, 'neigh_op_bnr_3')
// (7, 0, 'span12_vert_13')
// (7, 0, 'span4_vert_40')
// (7, 1, 'sp12_v_b_13')
// (7, 1, 'sp4_v_b_40')
// (7, 2, 'sp12_v_b_10')
// (7, 2, 'sp4_v_b_29')
// (7, 3, 'local_g2_1')
// (7, 3, 'lutff_2/in_3')
// (7, 3, 'lutff_7/in_0')
// (7, 3, 'neigh_op_top_3')
// (7, 3, 'sp12_v_b_9')
// (7, 3, 'sp4_v_b_16')
// (7, 4, 'local_g0_3')
// (7, 4, 'lutff_3/out')
// (7, 4, 'lutff_5/in_2')
// (7, 4, 'sp12_v_b_6')
// (7, 4, 'sp4_h_r_5')
// (7, 4, 'sp4_v_b_5')
// (7, 5, 'neigh_op_bot_3')
// (7, 5, 'sp12_v_b_5')
// (7, 6, 'sp12_v_b_2')
// (7, 7, 'sp12_v_b_1')
// (8, 3, 'local_g3_3')
// (8, 3, 'lutff_1/in_1')
// (8, 3, 'neigh_op_tnl_3')
// (8, 4, 'local_g0_0')
// (8, 4, 'lutff_4/in_2')
// (8, 4, 'lutff_5/in_1')
// (8, 4, 'neigh_op_lft_3')
// (8, 4, 'sp4_h_r_16')
// (8, 5, 'neigh_op_bnl_3')
// (9, 4, 'sp4_h_r_29')
// (10, 4, 'sp4_h_r_40')
// (11, 4, 'sp4_h_l_40')

wire n315;
// (6, 1, 'sp4_r_v_b_41')
// (6, 2, 'sp4_r_v_b_28')
// (6, 3, 'neigh_op_tnr_2')
// (6, 3, 'sp4_r_v_b_17')
// (6, 4, 'neigh_op_rgt_2')
// (6, 4, 'sp4_r_v_b_4')
// (6, 5, 'neigh_op_bnr_2')
// (7, 0, 'span4_vert_41')
// (7, 1, 'sp4_v_b_41')
// (7, 2, 'sp4_r_v_b_45')
// (7, 2, 'sp4_v_b_28')
// (7, 3, 'local_g0_1')
// (7, 3, 'local_g0_3')
// (7, 3, 'lutff_3/in_2')
// (7, 3, 'lutff_4/in_3')
// (7, 3, 'neigh_op_top_2')
// (7, 3, 'sp4_r_v_b_32')
// (7, 3, 'sp4_v_b_17')
// (7, 4, 'local_g0_2')
// (7, 4, 'lutff_2/out')
// (7, 4, 'lutff_5/in_1')
// (7, 4, 'sp4_r_v_b_21')
// (7, 4, 'sp4_v_b_4')
// (7, 5, 'neigh_op_bot_2')
// (7, 5, 'sp4_r_v_b_8')
// (8, 1, 'sp4_v_t_45')
// (8, 2, 'sp4_v_b_45')
// (8, 3, 'local_g2_2')
// (8, 3, 'local_g3_2')
// (8, 3, 'lutff_0/in_1')
// (8, 3, 'lutff_5/in_3')
// (8, 3, 'neigh_op_tnl_2')
// (8, 3, 'sp4_v_b_32')
// (8, 4, 'neigh_op_lft_2')
// (8, 4, 'sp4_v_b_21')
// (8, 5, 'neigh_op_bnl_2')
// (8, 5, 'sp4_v_b_8')

wire n316;
// (6, 2, 'neigh_op_tnr_0')
// (6, 3, 'neigh_op_rgt_0')
// (6, 4, 'neigh_op_bnr_0')
// (7, 2, 'local_g0_0')
// (7, 2, 'local_g1_0')
// (7, 2, 'lutff_4/in_1')
// (7, 2, 'lutff_7/in_1')
// (7, 2, 'neigh_op_top_0')
// (7, 3, 'lutff_0/out')
// (7, 4, 'neigh_op_bot_0')
// (8, 2, 'neigh_op_tnl_0')
// (8, 3, 'neigh_op_lft_0')
// (8, 4, 'neigh_op_bnl_0')

wire n317;
// (6, 2, 'neigh_op_tnr_1')
// (6, 3, 'neigh_op_rgt_1')
// (6, 4, 'neigh_op_bnr_1')
// (7, 0, 'span12_vert_6')
// (7, 1, 'sp12_v_b_6')
// (7, 2, 'local_g1_1')
// (7, 2, 'local_g2_5')
// (7, 2, 'lutff_2/in_3')
// (7, 2, 'lutff_5/in_3')
// (7, 2, 'neigh_op_top_1')
// (7, 2, 'sp12_v_b_5')
// (7, 3, 'lutff_1/out')
// (7, 3, 'sp12_v_b_2')
// (7, 4, 'neigh_op_bot_1')
// (7, 4, 'sp12_v_b_1')
// (8, 2, 'neigh_op_tnl_1')
// (8, 3, 'neigh_op_lft_1')
// (8, 4, 'neigh_op_bnl_1')

wire n318;
// (6, 2, 'neigh_op_tnr_2')
// (6, 3, 'neigh_op_rgt_2')
// (6, 4, 'neigh_op_bnr_2')
// (7, 2, 'local_g0_2')
// (7, 2, 'local_g1_2')
// (7, 2, 'lutff_4/in_3')
// (7, 2, 'lutff_7/in_3')
// (7, 2, 'neigh_op_top_2')
// (7, 3, 'local_g0_2')
// (7, 3, 'local_g1_2')
// (7, 3, 'lutff_1/in_2')
// (7, 3, 'lutff_2/out')
// (7, 3, 'lutff_6/in_2')
// (7, 4, 'neigh_op_bot_2')
// (8, 2, 'neigh_op_tnl_2')
// (8, 3, 'neigh_op_lft_2')
// (8, 4, 'neigh_op_bnl_2')

wire n319;
// (6, 2, 'neigh_op_tnr_3')
// (6, 3, 'neigh_op_rgt_3')
// (6, 4, 'neigh_op_bnr_3')
// (7, 2, 'neigh_op_top_3')
// (7, 3, 'local_g1_3')
// (7, 3, 'lutff_1/in_3')
// (7, 3, 'lutff_3/out')
// (7, 4, 'neigh_op_bot_3')
// (8, 2, 'neigh_op_tnl_3')
// (8, 3, 'neigh_op_lft_3')
// (8, 4, 'neigh_op_bnl_3')

wire n320;
// (6, 2, 'neigh_op_tnr_4')
// (6, 3, 'neigh_op_rgt_4')
// (6, 4, 'neigh_op_bnr_4')
// (7, 2, 'neigh_op_top_4')
// (7, 3, 'local_g1_4')
// (7, 3, 'lutff_4/out')
// (7, 3, 'lutff_6/in_3')
// (7, 4, 'neigh_op_bot_4')
// (8, 2, 'neigh_op_tnl_4')
// (8, 3, 'neigh_op_lft_4')
// (8, 4, 'neigh_op_bnl_4')

wire n321;
// (6, 2, 'neigh_op_tnr_5')
// (6, 2, 'sp4_r_v_b_39')
// (6, 3, 'neigh_op_rgt_5')
// (6, 3, 'sp4_r_v_b_26')
// (6, 4, 'neigh_op_bnr_5')
// (6, 4, 'sp4_r_v_b_15')
// (6, 5, 'sp4_r_v_b_2')
// (7, 1, 'sp4_v_t_39')
// (7, 2, 'local_g1_5')
// (7, 2, 'local_g2_7')
// (7, 2, 'lutff_0/in_3')
// (7, 2, 'lutff_3/in_3')
// (7, 2, 'lutff_6/in_0')
// (7, 2, 'neigh_op_top_5')
// (7, 2, 'sp4_v_b_39')
// (7, 3, 'lutff_5/out')
// (7, 3, 'sp4_v_b_26')
// (7, 4, 'neigh_op_bot_5')
// (7, 4, 'sp4_v_b_15')
// (7, 5, 'sp4_v_b_2')
// (8, 2, 'neigh_op_tnl_5')
// (8, 3, 'neigh_op_lft_5')
// (8, 4, 'neigh_op_bnl_5')

wire n322;
// (6, 3, 'neigh_op_tnr_0')
// (6, 4, 'neigh_op_rgt_0')
// (6, 5, 'neigh_op_bnr_0')
// (7, 3, 'neigh_op_top_0')
// (7, 4, 'local_g1_0')
// (7, 4, 'lutff_0/out')
// (7, 4, 'lutff_7/in_2')
// (7, 5, 'neigh_op_bot_0')
// (8, 3, 'local_g2_0')
// (8, 3, 'local_g3_0')
// (8, 3, 'lutff_2/in_1')
// (8, 3, 'lutff_3/in_3')
// (8, 3, 'neigh_op_tnl_0')
// (8, 4, 'neigh_op_lft_0')
// (8, 5, 'neigh_op_bnl_0')

wire n323;
// (6, 3, 'neigh_op_tnr_1')
// (6, 4, 'neigh_op_rgt_1')
// (6, 5, 'neigh_op_bnr_1')
// (7, 3, 'neigh_op_top_1')
// (7, 4, 'lutff_1/out')
// (7, 5, 'local_g1_1')
// (7, 5, 'lutff_6/in_2')
// (7, 5, 'neigh_op_bot_1')
// (8, 3, 'neigh_op_tnl_1')
// (8, 4, 'neigh_op_lft_1')
// (8, 5, 'neigh_op_bnl_1')

wire n324;
// (6, 3, 'neigh_op_tnr_4')
// (6, 4, 'neigh_op_rgt_4')
// (6, 5, 'neigh_op_bnr_4')
// (7, 0, 'span12_vert_15')
// (7, 1, 'sp12_v_b_15')
// (7, 2, 'sp12_v_b_12')
// (7, 3, 'local_g0_4')
// (7, 3, 'local_g2_3')
// (7, 3, 'lutff_3/in_0')
// (7, 3, 'lutff_4/in_0')
// (7, 3, 'neigh_op_top_4')
// (7, 3, 'sp12_v_b_11')
// (7, 4, 'lutff_4/out')
// (7, 4, 'sp12_v_b_8')
// (7, 5, 'neigh_op_bot_4')
// (7, 5, 'sp12_v_b_7')
// (7, 6, 'sp12_v_b_4')
// (7, 7, 'sp12_v_b_3')
// (7, 8, 'sp12_v_b_0')
// (8, 3, 'local_g2_4')
// (8, 3, 'local_g3_4')
// (8, 3, 'lutff_2/in_3')
// (8, 3, 'lutff_3/in_1')
// (8, 3, 'neigh_op_tnl_4')
// (8, 4, 'neigh_op_lft_4')
// (8, 5, 'neigh_op_bnl_4')

wire n325;
// (6, 3, 'neigh_op_tnr_5')
// (6, 4, 'neigh_op_rgt_5')
// (6, 4, 'sp12_h_r_1')
// (6, 4, 'sp4_h_r_0')
// (6, 5, 'neigh_op_bnr_5')
// (7, 3, 'local_g0_5')
// (7, 3, 'lutff_0/in_1')
// (7, 3, 'lutff_6/in_1')
// (7, 3, 'neigh_op_top_5')
// (7, 4, 'lutff_5/out')
// (7, 4, 'sp12_h_r_2')
// (7, 4, 'sp4_h_r_13')
// (7, 5, 'neigh_op_bot_5')
// (8, 3, 'local_g2_5')
// (8, 3, 'local_g3_5')
// (8, 3, 'lutff_1/in_2')
// (8, 3, 'lutff_7/in_3')
// (8, 3, 'neigh_op_tnl_5')
// (8, 4, 'local_g2_0')
// (8, 4, 'lutff_7/in_3')
// (8, 4, 'neigh_op_lft_5')
// (8, 4, 'sp12_h_r_5')
// (8, 4, 'sp4_h_r_24')
// (8, 5, 'neigh_op_bnl_5')
// (9, 4, 'sp12_h_r_6')
// (9, 4, 'sp4_h_r_37')
// (10, 4, 'sp12_h_r_9')
// (10, 4, 'sp4_h_l_37')
// (11, 4, 'sp12_h_r_10')
// (12, 4, 'sp12_h_r_13')
// (13, 4, 'span12_horz_13')

wire n326;
// (6, 3, 'neigh_op_tnr_6')
// (6, 4, 'neigh_op_rgt_6')
// (6, 5, 'neigh_op_bnr_6')
// (7, 3, 'local_g0_6')
// (7, 3, 'local_g1_6')
// (7, 3, 'lutff_0/in_2')
// (7, 3, 'lutff_5/in_2')
// (7, 3, 'neigh_op_top_6')
// (7, 4, 'local_g2_6')
// (7, 4, 'lutff_1/in_1')
// (7, 4, 'lutff_6/out')
// (7, 5, 'neigh_op_bot_6')
// (8, 3, 'neigh_op_tnl_6')
// (8, 4, 'neigh_op_lft_6')
// (8, 5, 'neigh_op_bnl_6')

wire n327;
// (6, 3, 'sp4_r_v_b_36')
// (6, 4, 'neigh_op_tnr_6')
// (6, 4, 'sp4_r_v_b_25')
// (6, 5, 'neigh_op_rgt_6')
// (6, 5, 'sp4_r_v_b_12')
// (6, 6, 'neigh_op_bnr_6')
// (6, 6, 'sp4_r_v_b_1')
// (7, 2, 'sp4_v_t_36')
// (7, 3, 'sp4_v_b_36')
// (7, 4, 'neigh_op_top_6')
// (7, 4, 'sp4_v_b_25')
// (7, 5, 'lutff_6/out')
// (7, 5, 'sp4_v_b_12')
// (7, 6, 'local_g0_1')
// (7, 6, 'lutff_0/in_1')
// (7, 6, 'neigh_op_bot_6')
// (7, 6, 'sp4_v_b_1')
// (8, 4, 'neigh_op_tnl_6')
// (8, 5, 'neigh_op_lft_6')
// (8, 6, 'neigh_op_bnl_6')

wire n328;
// (6, 4, 'neigh_op_tnr_0')
// (6, 5, 'neigh_op_rgt_0')
// (6, 6, 'neigh_op_bnr_0')
// (7, 4, 'neigh_op_top_0')
// (7, 5, 'local_g1_0')
// (7, 5, 'lutff_0/out')
// (7, 5, 'lutff_3/in_2')
// (7, 6, 'neigh_op_bot_0')
// (8, 4, 'neigh_op_tnl_0')
// (8, 5, 'neigh_op_lft_0')
// (8, 6, 'neigh_op_bnl_0')

wire n329;
// (6, 4, 'neigh_op_tnr_1')
// (6, 5, 'neigh_op_rgt_1')
// (6, 6, 'neigh_op_bnr_1')
// (7, 3, 'sp4_r_v_b_43')
// (7, 4, 'local_g1_6')
// (7, 4, 'lutff_3/in_2')
// (7, 4, 'lutff_6/in_3')
// (7, 4, 'neigh_op_top_1')
// (7, 4, 'sp4_r_v_b_30')
// (7, 5, 'lutff_1/out')
// (7, 5, 'sp4_r_v_b_19')
// (7, 6, 'neigh_op_bot_1')
// (7, 6, 'sp4_r_v_b_6')
// (8, 2, 'sp4_v_t_43')
// (8, 3, 'sp4_v_b_43')
// (8, 4, 'neigh_op_tnl_1')
// (8, 4, 'sp4_v_b_30')
// (8, 5, 'neigh_op_lft_1')
// (8, 5, 'sp4_v_b_19')
// (8, 6, 'neigh_op_bnl_1')
// (8, 6, 'sp4_v_b_6')

wire n330;
// (6, 4, 'neigh_op_tnr_2')
// (6, 5, 'neigh_op_rgt_2')
// (6, 6, 'neigh_op_bnr_2')
// (7, 4, 'neigh_op_top_2')
// (7, 5, 'local_g1_2')
// (7, 5, 'lutff_0/in_3')
// (7, 5, 'lutff_2/out')
// (7, 6, 'neigh_op_bot_2')
// (8, 4, 'neigh_op_tnl_2')
// (8, 5, 'neigh_op_lft_2')
// (8, 6, 'neigh_op_bnl_2')

wire n331;
// (6, 4, 'neigh_op_tnr_3')
// (6, 5, 'neigh_op_rgt_3')
// (6, 6, 'neigh_op_bnr_3')
// (7, 4, 'neigh_op_top_3')
// (7, 5, 'lutff_3/out')
// (7, 6, 'local_g0_3')
// (7, 6, 'lutff_1/in_2')
// (7, 6, 'neigh_op_bot_3')
// (8, 4, 'neigh_op_tnl_3')
// (8, 5, 'neigh_op_lft_3')
// (8, 6, 'neigh_op_bnl_3')

wire n332;
// (6, 4, 'neigh_op_tnr_5')
// (6, 5, 'neigh_op_rgt_5')
// (6, 6, 'neigh_op_bnr_5')
// (7, 4, 'neigh_op_top_5')
// (7, 5, 'lutff_5/out')
// (7, 6, 'neigh_op_bot_5')
// (8, 4, 'neigh_op_tnl_5')
// (8, 5, 'local_g0_5')
// (8, 5, 'lutff_2/in_1')
// (8, 5, 'neigh_op_lft_5')
// (8, 6, 'neigh_op_bnl_5')

reg n333 = 0;
// (6, 4, 'sp4_r_v_b_38')
// (6, 5, 'local_g0_3')
// (6, 5, 'lutff_0/in_3')
// (6, 5, 'sp4_r_v_b_27')
// (6, 6, 'sp4_r_v_b_14')
// (6, 7, 'sp4_r_v_b_3')
// (7, 3, 'sp4_v_t_38')
// (7, 4, 'sp4_v_b_38')
// (7, 5, 'sp4_v_b_27')
// (7, 6, 'sp4_v_b_14')
// (7, 7, 'sp4_h_r_3')
// (7, 7, 'sp4_v_b_3')
// (8, 7, 'sp4_h_r_14')
// (9, 7, 'sp4_h_r_27')
// (10, 7, 'neigh_op_tnr_3')
// (10, 7, 'sp4_h_r_38')
// (10, 8, 'neigh_op_rgt_3')
// (10, 8, 'sp4_r_v_b_38')
// (10, 9, 'neigh_op_bnr_3')
// (10, 9, 'sp4_r_v_b_27')
// (10, 10, 'sp4_r_v_b_14')
// (10, 11, 'sp4_r_v_b_3')
// (11, 7, 'neigh_op_top_3')
// (11, 7, 'sp4_h_l_38')
// (11, 7, 'sp4_v_t_38')
// (11, 8, 'local_g1_3')
// (11, 8, 'lutff_3/out')
// (11, 8, 'lutff_4/in_0')
// (11, 8, 'sp4_v_b_38')
// (11, 9, 'neigh_op_bot_3')
// (11, 9, 'sp4_v_b_27')
// (11, 10, 'sp4_v_b_14')
// (11, 11, 'sp4_v_b_3')
// (12, 7, 'neigh_op_tnl_3')
// (12, 8, 'neigh_op_lft_3')
// (12, 9, 'neigh_op_bnl_3')

wire n334;
// (6, 5, 'neigh_op_tnr_2')
// (6, 6, 'neigh_op_rgt_2')
// (6, 7, 'neigh_op_bnr_2')
// (7, 5, 'neigh_op_top_2')
// (7, 6, 'local_g0_2')
// (7, 6, 'lutff_0/in_2')
// (7, 6, 'lutff_2/out')
// (7, 7, 'neigh_op_bot_2')
// (8, 5, 'neigh_op_tnl_2')
// (8, 6, 'neigh_op_lft_2')
// (8, 7, 'neigh_op_bnl_2')

wire n335;
// (6, 5, 'neigh_op_tnr_3')
// (6, 6, 'neigh_op_rgt_3')
// (6, 7, 'neigh_op_bnr_3')
// (7, 5, 'neigh_op_top_3')
// (7, 6, 'local_g1_3')
// (7, 6, 'lutff_3/out')
// (7, 6, 'lutff_6/in_2')
// (7, 7, 'neigh_op_bot_3')
// (8, 5, 'local_g3_3')
// (8, 5, 'lutff_2/in_0')
// (8, 5, 'neigh_op_tnl_3')
// (8, 6, 'neigh_op_lft_3')
// (8, 7, 'neigh_op_bnl_3')

wire n336;
// (6, 5, 'neigh_op_tnr_4')
// (6, 6, 'neigh_op_rgt_4')
// (6, 7, 'neigh_op_bnr_4')
// (7, 5, 'neigh_op_top_4')
// (7, 6, 'local_g0_4')
// (7, 6, 'lutff_2/in_2')
// (7, 6, 'lutff_4/out')
// (7, 7, 'neigh_op_bot_4')
// (8, 5, 'neigh_op_tnl_4')
// (8, 6, 'neigh_op_lft_4')
// (8, 7, 'neigh_op_bnl_4')

wire n337;
// (6, 5, 'neigh_op_tnr_6')
// (6, 6, 'neigh_op_rgt_6')
// (6, 7, 'neigh_op_bnr_6')
// (7, 5, 'neigh_op_top_6')
// (7, 6, 'local_g1_6')
// (7, 6, 'lutff_5/in_2')
// (7, 6, 'lutff_6/out')
// (7, 7, 'neigh_op_bot_6')
// (8, 5, 'neigh_op_tnl_6')
// (8, 6, 'neigh_op_lft_6')
// (8, 7, 'neigh_op_bnl_6')

reg n338 = 0;
// (6, 5, 'neigh_op_tnr_7')
// (6, 6, 'neigh_op_rgt_7')
// (6, 7, 'neigh_op_bnr_7')
// (7, 5, 'local_g1_7')
// (7, 5, 'lutff_1/in_1')
// (7, 5, 'neigh_op_top_7')
// (7, 6, 'lutff_7/out')
// (7, 7, 'neigh_op_bot_7')
// (8, 5, 'neigh_op_tnl_7')
// (8, 6, 'neigh_op_lft_7')
// (8, 7, 'neigh_op_bnl_7')

wire n339;
// (6, 5, 'sp4_r_v_b_44')
// (6, 6, 'neigh_op_tnr_2')
// (6, 6, 'sp4_r_v_b_33')
// (6, 7, 'neigh_op_rgt_2')
// (6, 7, 'sp4_r_v_b_20')
// (6, 8, 'neigh_op_bnr_2')
// (6, 8, 'sp4_r_v_b_9')
// (7, 4, 'sp4_v_t_44')
// (7, 5, 'sp4_v_b_44')
// (7, 6, 'neigh_op_top_2')
// (7, 6, 'sp4_v_b_33')
// (7, 7, 'lutff_2/out')
// (7, 7, 'sp4_r_v_b_37')
// (7, 7, 'sp4_v_b_20')
// (7, 8, 'local_g1_0')
// (7, 8, 'local_g1_1')
// (7, 8, 'lutff_0/in_2')
// (7, 8, 'lutff_6/in_3')
// (7, 8, 'lutff_7/in_2')
// (7, 8, 'neigh_op_bot_2')
// (7, 8, 'sp4_r_v_b_24')
// (7, 8, 'sp4_v_b_9')
// (7, 9, 'sp4_r_v_b_13')
// (7, 10, 'sp4_r_v_b_0')
// (8, 6, 'local_g2_2')
// (8, 6, 'lutff_2/in_0')
// (8, 6, 'lutff_4/in_0')
// (8, 6, 'lutff_5/in_3')
// (8, 6, 'lutff_6/in_0')
// (8, 6, 'neigh_op_tnl_2')
// (8, 6, 'sp4_v_t_37')
// (8, 7, 'local_g2_5')
// (8, 7, 'lutff_1/in_0')
// (8, 7, 'neigh_op_lft_2')
// (8, 7, 'sp4_v_b_37')
// (8, 8, 'neigh_op_bnl_2')
// (8, 8, 'sp4_v_b_24')
// (8, 9, 'sp4_v_b_13')
// (8, 10, 'sp4_v_b_0')

reg n340 = 0;
// (6, 5, 'sp4_r_v_b_46')
// (6, 6, 'local_g0_0')
// (6, 6, 'lutff_6/in_0')
// (6, 6, 'sp4_r_v_b_35')
// (6, 7, 'sp4_r_v_b_22')
// (6, 8, 'sp4_r_v_b_11')
// (6, 9, 'sp4_r_v_b_40')
// (6, 10, 'sp4_r_v_b_29')
// (6, 11, 'sp4_r_v_b_16')
// (6, 12, 'sp4_r_v_b_5')
// (6, 13, 'sp4_r_v_b_36')
// (6, 14, 'sp4_r_v_b_25')
// (6, 15, 'sp4_r_v_b_12')
// (6, 16, 'sp4_r_v_b_1')
// (7, 4, 'sp4_v_t_46')
// (7, 5, 'sp4_v_b_46')
// (7, 6, 'sp4_v_b_35')
// (7, 7, 'sp4_v_b_22')
// (7, 8, 'sp4_h_r_11')
// (7, 8, 'sp4_v_b_11')
// (7, 8, 'sp4_v_t_40')
// (7, 9, 'sp4_v_b_40')
// (7, 10, 'local_g3_5')
// (7, 10, 'lutff_0/in_2')
// (7, 10, 'sp4_v_b_29')
// (7, 11, 'sp4_v_b_16')
// (7, 12, 'sp4_v_b_5')
// (7, 12, 'sp4_v_t_36')
// (7, 13, 'local_g2_4')
// (7, 13, 'lutff_0/in_2')
// (7, 13, 'sp4_v_b_36')
// (7, 14, 'sp4_v_b_25')
// (7, 15, 'sp4_v_b_12')
// (7, 16, 'sp4_v_b_1')
// (8, 8, 'sp4_h_r_22')
// (8, 9, 'sp4_r_v_b_43')
// (8, 10, 'sp4_r_v_b_30')
// (8, 11, 'sp4_r_v_b_19')
// (8, 12, 'sp4_r_v_b_6')
// (8, 13, 'sp4_r_v_b_43')
// (8, 14, 'sp4_r_v_b_30')
// (8, 15, 'sp4_r_v_b_19')
// (8, 16, 'sp4_r_v_b_6')
// (9, 8, 'sp4_h_r_0')
// (9, 8, 'sp4_h_r_35')
// (9, 8, 'sp4_v_t_43')
// (9, 9, 'sp4_v_b_43')
// (9, 10, 'sp4_v_b_30')
// (9, 11, 'sp4_v_b_19')
// (9, 12, 'sp4_v_b_6')
// (9, 12, 'sp4_v_t_43')
// (9, 13, 'local_g2_3')
// (9, 13, 'lutff_7/in_0')
// (9, 13, 'sp4_v_b_43')
// (9, 14, 'sp4_v_b_30')
// (9, 15, 'sp4_v_b_19')
// (9, 16, 'sp4_v_b_6')
// (10, 7, 'neigh_op_tnr_4')
// (10, 8, 'neigh_op_rgt_4')
// (10, 8, 'sp4_h_r_13')
// (10, 8, 'sp4_h_r_46')
// (10, 9, 'neigh_op_bnr_4')
// (11, 7, 'neigh_op_top_4')
// (11, 8, 'lutff_4/out')
// (11, 8, 'sp4_h_l_46')
// (11, 8, 'sp4_h_r_24')
// (11, 8, 'sp4_h_r_8')
// (11, 9, 'neigh_op_bot_4')
// (12, 7, 'neigh_op_tnl_4')
// (12, 8, 'neigh_op_lft_4')
// (12, 8, 'sp4_h_r_21')
// (12, 8, 'sp4_h_r_37')
// (12, 9, 'neigh_op_bnl_4')
// (13, 8, 'span4_horz_21')
// (13, 8, 'span4_horz_37')

wire n341;
// (6, 5, 'sp4_r_v_b_47')
// (6, 6, 'sp4_r_v_b_34')
// (6, 7, 'neigh_op_tnr_5')
// (6, 7, 'sp4_r_v_b_23')
// (6, 8, 'neigh_op_rgt_5')
// (6, 8, 'sp4_r_v_b_10')
// (6, 9, 'neigh_op_bnr_5')
// (7, 4, 'sp4_v_t_47')
// (7, 5, 'sp4_v_b_47')
// (7, 6, 'sp4_v_b_34')
// (7, 7, 'local_g1_7')
// (7, 7, 'lutff_2/in_2')
// (7, 7, 'neigh_op_top_5')
// (7, 7, 'sp4_v_b_23')
// (7, 8, 'lutff_5/out')
// (7, 8, 'sp4_v_b_10')
// (7, 9, 'neigh_op_bot_5')
// (8, 7, 'neigh_op_tnl_5')
// (8, 8, 'neigh_op_lft_5')
// (8, 9, 'neigh_op_bnl_5')

wire n342;
// (6, 6, 'neigh_op_tnr_0')
// (6, 7, 'neigh_op_rgt_0')
// (6, 8, 'neigh_op_bnr_0')
// (7, 6, 'neigh_op_top_0')
// (7, 7, 'local_g1_0')
// (7, 7, 'local_g2_0')
// (7, 7, 'lutff_0/out')
// (7, 7, 'lutff_2/in_3')
// (7, 7, 'lutff_7/in_1')
// (7, 8, 'neigh_op_bot_0')
// (8, 6, 'neigh_op_tnl_0')
// (8, 7, 'neigh_op_lft_0')
// (8, 8, 'neigh_op_bnl_0')

wire n343;
// (6, 6, 'neigh_op_tnr_1')
// (6, 7, 'neigh_op_rgt_1')
// (6, 8, 'neigh_op_bnr_1')
// (7, 6, 'neigh_op_top_1')
// (7, 7, 'local_g3_1')
// (7, 7, 'lutff_1/out')
// (7, 7, 'lutff_7/in_3')
// (7, 8, 'neigh_op_bot_1')
// (8, 6, 'neigh_op_tnl_1')
// (8, 7, 'neigh_op_lft_1')
// (8, 8, 'neigh_op_bnl_1')

wire n344;
// (6, 6, 'neigh_op_tnr_3')
// (6, 7, 'neigh_op_rgt_3')
// (6, 8, 'neigh_op_bnr_3')
// (7, 6, 'neigh_op_top_3')
// (7, 7, 'local_g2_3')
// (7, 7, 'lutff_3/out')
// (7, 7, 'lutff_5/in_2')
// (7, 7, 'lutff_7/in_2')
// (7, 8, 'neigh_op_bot_3')
// (8, 6, 'neigh_op_tnl_3')
// (8, 7, 'neigh_op_lft_3')
// (8, 8, 'neigh_op_bnl_3')

wire n345;
// (6, 6, 'neigh_op_tnr_4')
// (6, 7, 'neigh_op_rgt_4')
// (6, 8, 'neigh_op_bnr_4')
// (7, 6, 'neigh_op_top_4')
// (7, 7, 'local_g2_4')
// (7, 7, 'lutff_4/out')
// (7, 7, 'lutff_5/in_3')
// (7, 8, 'neigh_op_bot_4')
// (8, 6, 'neigh_op_tnl_4')
// (8, 7, 'neigh_op_lft_4')
// (8, 8, 'neigh_op_bnl_4')

wire n346;
// (6, 6, 'neigh_op_tnr_5')
// (6, 7, 'neigh_op_rgt_5')
// (6, 8, 'neigh_op_bnr_5')
// (7, 0, 'span12_vert_22')
// (7, 1, 'sp12_v_b_22')
// (7, 2, 'sp12_v_b_21')
// (7, 3, 'sp12_v_b_18')
// (7, 4, 'sp12_v_b_17')
// (7, 5, 'sp12_v_b_14')
// (7, 6, 'neigh_op_top_5')
// (7, 6, 'sp12_v_b_13')
// (7, 6, 'sp4_r_v_b_38')
// (7, 7, 'lutff_5/out')
// (7, 7, 'sp12_v_b_10')
// (7, 7, 'sp4_r_v_b_27')
// (7, 8, 'local_g2_1')
// (7, 8, 'local_g3_1')
// (7, 8, 'lutff_0/in_3')
// (7, 8, 'lutff_6/in_1')
// (7, 8, 'lutff_7/in_1')
// (7, 8, 'neigh_op_bot_5')
// (7, 8, 'sp12_v_b_9')
// (7, 8, 'sp4_r_v_b_14')
// (7, 9, 'sp12_v_b_6')
// (7, 9, 'sp4_r_v_b_3')
// (7, 10, 'sp12_v_b_5')
// (7, 11, 'sp12_v_b_2')
// (7, 12, 'sp12_v_b_1')
// (8, 5, 'sp4_v_t_38')
// (8, 6, 'local_g2_5')
// (8, 6, 'local_g3_5')
// (8, 6, 'lutff_2/in_3')
// (8, 6, 'lutff_4/in_2')
// (8, 6, 'lutff_5/in_2')
// (8, 6, 'lutff_6/in_2')
// (8, 6, 'neigh_op_tnl_5')
// (8, 6, 'sp4_v_b_38')
// (8, 7, 'local_g3_3')
// (8, 7, 'lutff_1/in_1')
// (8, 7, 'neigh_op_lft_5')
// (8, 7, 'sp4_v_b_27')
// (8, 8, 'neigh_op_bnl_5')
// (8, 8, 'sp4_v_b_14')
// (8, 9, 'sp4_v_b_3')

wire n347;
// (6, 6, 'neigh_op_tnr_6')
// (6, 7, 'neigh_op_rgt_6')
// (6, 8, 'neigh_op_bnr_6')
// (7, 6, 'neigh_op_top_6')
// (7, 7, 'local_g1_6')
// (7, 7, 'lutff_0/in_1')
// (7, 7, 'lutff_1/in_2')
// (7, 7, 'lutff_6/out')
// (7, 8, 'neigh_op_bot_6')
// (8, 6, 'neigh_op_tnl_6')
// (8, 7, 'local_g1_6')
// (8, 7, 'lutff_4/in_1')
// (8, 7, 'lutff_6/in_3')
// (8, 7, 'neigh_op_lft_6')
// (8, 8, 'neigh_op_bnl_6')

wire n348;
// (6, 7, 'neigh_op_tnr_0')
// (6, 8, 'neigh_op_rgt_0')
// (6, 9, 'neigh_op_bnr_0')
// (7, 7, 'neigh_op_top_0')
// (7, 8, 'local_g2_0')
// (7, 8, 'local_g3_0')
// (7, 8, 'lutff_0/out')
// (7, 8, 'lutff_1/in_0')
// (7, 8, 'lutff_2/in_0')
// (7, 9, 'neigh_op_bot_0')
// (8, 7, 'neigh_op_tnl_0')
// (8, 8, 'neigh_op_lft_0')
// (8, 9, 'neigh_op_bnl_0')

wire n349;
// (6, 7, 'neigh_op_tnr_2')
// (6, 8, 'neigh_op_rgt_2')
// (6, 9, 'neigh_op_bnr_2')
// (7, 7, 'neigh_op_top_2')
// (7, 8, 'lutff_2/out')
// (7, 9, 'neigh_op_bot_2')
// (8, 7, 'local_g2_2')
// (8, 7, 'lutff_2/in_2')
// (8, 7, 'neigh_op_tnl_2')
// (8, 8, 'local_g0_2')
// (8, 8, 'lutff_1/in_3')
// (8, 8, 'neigh_op_lft_2')
// (8, 9, 'neigh_op_bnl_2')

wire n350;
// (6, 7, 'neigh_op_tnr_3')
// (6, 8, 'neigh_op_rgt_3')
// (6, 9, 'neigh_op_bnr_3')
// (7, 7, 'neigh_op_top_3')
// (7, 8, 'lutff_3/out')
// (7, 9, 'neigh_op_bot_3')
// (8, 7, 'neigh_op_tnl_3')
// (8, 8, 'local_g1_3')
// (8, 8, 'lutff_5/in_3')
// (8, 8, 'neigh_op_lft_3')
// (8, 9, 'neigh_op_bnl_3')

wire n351;
// (6, 7, 'neigh_op_tnr_6')
// (6, 8, 'neigh_op_rgt_6')
// (6, 9, 'neigh_op_bnr_6')
// (7, 7, 'neigh_op_top_6')
// (7, 8, 'local_g1_6')
// (7, 8, 'lutff_3/in_0')
// (7, 8, 'lutff_4/in_1')
// (7, 8, 'lutff_6/out')
// (7, 9, 'neigh_op_bot_6')
// (8, 7, 'neigh_op_tnl_6')
// (8, 8, 'neigh_op_lft_6')
// (8, 9, 'neigh_op_bnl_6')

wire n352;
// (6, 7, 'neigh_op_tnr_7')
// (6, 8, 'neigh_op_rgt_7')
// (6, 9, 'neigh_op_bnr_7')
// (7, 7, 'neigh_op_top_7')
// (7, 8, 'local_g0_7')
// (7, 8, 'local_g1_7')
// (7, 8, 'lutff_1/in_2')
// (7, 8, 'lutff_2/in_2')
// (7, 8, 'lutff_3/in_2')
// (7, 8, 'lutff_4/in_2')
// (7, 8, 'lutff_7/out')
// (7, 9, 'neigh_op_bot_7')
// (8, 7, 'neigh_op_tnl_7')
// (8, 8, 'neigh_op_lft_7')
// (8, 9, 'neigh_op_bnl_7')

wire n353;
// (6, 8, 'neigh_op_tnr_0')
// (6, 9, 'local_g2_0')
// (6, 9, 'lutff_3/in_1')
// (6, 9, 'lutff_7/in_1')
// (6, 9, 'neigh_op_rgt_0')
// (6, 10, 'neigh_op_bnr_0')
// (7, 8, 'neigh_op_top_0')
// (7, 9, 'lutff_0/out')
// (7, 10, 'neigh_op_bot_0')
// (8, 8, 'neigh_op_tnl_0')
// (8, 9, 'neigh_op_lft_0')
// (8, 10, 'neigh_op_bnl_0')

reg n354 = 0;
// (6, 8, 'neigh_op_tnr_1')
// (6, 9, 'neigh_op_rgt_1')
// (6, 10, 'neigh_op_bnr_1')
// (7, 8, 'neigh_op_top_1')
// (7, 9, 'local_g0_1')
// (7, 9, 'lutff_1/out')
// (7, 9, 'lutff_5/in_0')
// (7, 10, 'neigh_op_bot_1')
// (8, 8, 'neigh_op_tnl_1')
// (8, 9, 'neigh_op_lft_1')
// (8, 10, 'neigh_op_bnl_1')

reg n355 = 0;
// (6, 8, 'neigh_op_tnr_2')
// (6, 9, 'neigh_op_rgt_2')
// (6, 10, 'neigh_op_bnr_2')
// (7, 8, 'neigh_op_top_2')
// (7, 9, 'local_g1_2')
// (7, 9, 'lutff_1/in_0')
// (7, 9, 'lutff_2/out')
// (7, 10, 'neigh_op_bot_2')
// (8, 8, 'neigh_op_tnl_2')
// (8, 9, 'neigh_op_lft_2')
// (8, 10, 'neigh_op_bnl_2')

reg n356 = 0;
// (6, 8, 'neigh_op_tnr_4')
// (6, 9, 'neigh_op_rgt_4')
// (6, 10, 'neigh_op_bnr_4')
// (7, 8, 'neigh_op_top_4')
// (7, 9, 'local_g0_4')
// (7, 9, 'lutff_4/out')
// (7, 9, 'lutff_6/in_0')
// (7, 10, 'neigh_op_bot_4')
// (8, 8, 'neigh_op_tnl_4')
// (8, 9, 'neigh_op_lft_4')
// (8, 10, 'neigh_op_bnl_4')

reg n357 = 0;
// (6, 8, 'neigh_op_tnr_5')
// (6, 9, 'neigh_op_rgt_5')
// (6, 10, 'neigh_op_bnr_5')
// (7, 8, 'neigh_op_top_5')
// (7, 9, 'local_g0_5')
// (7, 9, 'lutff_3/in_0')
// (7, 9, 'lutff_5/out')
// (7, 10, 'neigh_op_bot_5')
// (8, 8, 'neigh_op_tnl_5')
// (8, 9, 'neigh_op_lft_5')
// (8, 10, 'neigh_op_bnl_5')

reg n358 = 0;
// (6, 8, 'neigh_op_tnr_6')
// (6, 9, 'neigh_op_rgt_6')
// (6, 10, 'neigh_op_bnr_6')
// (7, 8, 'neigh_op_top_6')
// (7, 8, 'sp4_r_v_b_40')
// (7, 9, 'lutff_6/out')
// (7, 9, 'sp4_r_v_b_29')
// (7, 10, 'neigh_op_bot_6')
// (7, 10, 'sp4_r_v_b_16')
// (7, 11, 'sp4_r_v_b_5')
// (8, 7, 'sp4_h_r_10')
// (8, 7, 'sp4_v_t_40')
// (8, 8, 'neigh_op_tnl_6')
// (8, 8, 'sp4_v_b_40')
// (8, 9, 'neigh_op_lft_6')
// (8, 9, 'sp4_v_b_29')
// (8, 10, 'neigh_op_bnl_6')
// (8, 10, 'sp4_v_b_16')
// (8, 11, 'sp4_v_b_5')
// (9, 7, 'sp4_h_r_23')
// (10, 7, 'sp4_h_r_34')
// (11, 7, 'local_g3_7')
// (11, 7, 'lutff_0/in_0')
// (11, 7, 'sp4_h_r_47')
// (12, 7, 'sp4_h_l_47')

wire n359;
// (6, 8, 'sp4_r_v_b_39')
// (6, 9, 'local_g0_2')
// (6, 9, 'local_g3_2')
// (6, 9, 'lutff_1/in_2')
// (6, 9, 'lutff_5/in_3')
// (6, 9, 'sp4_r_v_b_26')
// (6, 9, 'sp4_r_v_b_42')
// (6, 10, 'neigh_op_tnr_1')
// (6, 10, 'sp4_r_v_b_15')
// (6, 10, 'sp4_r_v_b_31')
// (6, 11, 'neigh_op_rgt_1')
// (6, 11, 'sp4_r_v_b_18')
// (6, 11, 'sp4_r_v_b_2')
// (6, 12, 'neigh_op_bnr_1')
// (6, 12, 'sp4_r_v_b_7')
// (7, 7, 'sp4_v_t_39')
// (7, 8, 'sp4_v_b_39')
// (7, 8, 'sp4_v_t_42')
// (7, 9, 'sp4_v_b_26')
// (7, 9, 'sp4_v_b_42')
// (7, 10, 'neigh_op_top_1')
// (7, 10, 'sp4_v_b_15')
// (7, 10, 'sp4_v_b_31')
// (7, 11, 'lutff_1/out')
// (7, 11, 'sp4_v_b_18')
// (7, 11, 'sp4_v_b_2')
// (7, 12, 'neigh_op_bot_1')
// (7, 12, 'sp4_v_b_7')
// (8, 10, 'neigh_op_tnl_1')
// (8, 11, 'neigh_op_lft_1')
// (8, 12, 'neigh_op_bnl_1')

wire n360;
// (6, 9, 'neigh_op_tnr_1')
// (6, 10, 'neigh_op_rgt_1')
// (6, 11, 'local_g0_1')
// (6, 11, 'lutff_0/in_1')
// (6, 11, 'lutff_4/in_1')
// (6, 11, 'neigh_op_bnr_1')
// (7, 9, 'neigh_op_top_1')
// (7, 10, 'lutff_1/out')
// (7, 11, 'neigh_op_bot_1')
// (8, 9, 'neigh_op_tnl_1')
// (8, 10, 'neigh_op_lft_1')
// (8, 11, 'neigh_op_bnl_1')

wire n361;
// (6, 9, 'neigh_op_tnr_2')
// (6, 10, 'neigh_op_rgt_2')
// (6, 11, 'neigh_op_bnr_2')
// (7, 9, 'neigh_op_top_2')
// (7, 10, 'local_g1_2')
// (7, 10, 'lutff_2/out')
// (7, 10, 'lutff_4/in_3')
// (7, 11, 'neigh_op_bot_2')
// (8, 9, 'neigh_op_tnl_2')
// (8, 10, 'neigh_op_lft_2')
// (8, 11, 'neigh_op_bnl_2')

wire n362;
// (6, 9, 'neigh_op_tnr_3')
// (6, 10, 'neigh_op_rgt_3')
// (6, 11, 'neigh_op_bnr_3')
// (7, 9, 'neigh_op_top_3')
// (7, 10, 'local_g0_3')
// (7, 10, 'lutff_2/in_3')
// (7, 10, 'lutff_3/out')
// (7, 11, 'neigh_op_bot_3')
// (8, 9, 'neigh_op_tnl_3')
// (8, 10, 'neigh_op_lft_3')
// (8, 11, 'neigh_op_bnl_3')

reg n363 = 0;
// (6, 9, 'neigh_op_tnr_5')
// (6, 10, 'local_g2_5')
// (6, 10, 'lutff_1/in_0')
// (6, 10, 'neigh_op_rgt_5')
// (6, 11, 'neigh_op_bnr_5')
// (7, 9, 'neigh_op_top_5')
// (7, 10, 'lutff_5/out')
// (7, 11, 'neigh_op_bot_5')
// (8, 9, 'neigh_op_tnl_5')
// (8, 10, 'neigh_op_lft_5')
// (8, 11, 'neigh_op_bnl_5')

reg n364 = 0;
// (6, 9, 'neigh_op_tnr_7')
// (6, 10, 'neigh_op_rgt_7')
// (6, 11, 'neigh_op_bnr_7')
// (7, 9, 'neigh_op_top_7')
// (7, 10, 'lutff_7/out')
// (7, 11, 'local_g0_7')
// (7, 11, 'lutff_5/in_0')
// (7, 11, 'neigh_op_bot_7')
// (8, 9, 'neigh_op_tnl_7')
// (8, 10, 'neigh_op_lft_7')
// (8, 11, 'neigh_op_bnl_7')

reg n365 = 0;
// (6, 9, 'sp4_r_v_b_43')
// (6, 10, 'sp4_r_v_b_30')
// (6, 11, 'neigh_op_tnr_6')
// (6, 11, 'sp4_r_v_b_19')
// (6, 12, 'neigh_op_rgt_6')
// (6, 12, 'sp4_r_v_b_6')
// (6, 13, 'neigh_op_bnr_6')
// (7, 6, 'sp12_v_t_23')
// (7, 7, 'sp12_v_b_23')
// (7, 8, 'sp12_v_b_20')
// (7, 8, 'sp4_v_t_43')
// (7, 9, 'sp12_v_b_19')
// (7, 9, 'sp4_v_b_43')
// (7, 10, 'local_g2_0')
// (7, 10, 'local_g3_6')
// (7, 10, 'lutff_2/in_0')
// (7, 10, 'lutff_5/in_0')
// (7, 10, 'lutff_7/in_0')
// (7, 10, 'sp12_v_b_16')
// (7, 10, 'sp4_v_b_30')
// (7, 11, 'neigh_op_top_6')
// (7, 11, 'sp12_v_b_15')
// (7, 11, 'sp4_v_b_19')
// (7, 12, 'local_g0_6')
// (7, 12, 'lutff_2/in_0')
// (7, 12, 'lutff_6/out')
// (7, 12, 'sp12_v_b_12')
// (7, 12, 'sp4_v_b_6')
// (7, 13, 'neigh_op_bot_6')
// (7, 13, 'sp12_v_b_11')
// (7, 14, 'sp12_v_b_8')
// (7, 15, 'sp12_v_b_7')
// (7, 16, 'sp12_v_b_4')
// (7, 17, 'span12_vert_3')
// (8, 11, 'neigh_op_tnl_6')
// (8, 12, 'neigh_op_lft_6')
// (8, 13, 'neigh_op_bnl_6')

wire n366;
// (6, 10, 'neigh_op_tnr_0')
// (6, 11, 'local_g2_0')
// (6, 11, 'lutff_1/in_1')
// (6, 11, 'neigh_op_rgt_0')
// (6, 12, 'local_g0_0')
// (6, 12, 'lutff_5/in_1')
// (6, 12, 'neigh_op_bnr_0')
// (7, 10, 'neigh_op_top_0')
// (7, 11, 'lutff_0/out')
// (7, 12, 'neigh_op_bot_0')
// (8, 10, 'neigh_op_tnl_0')
// (8, 11, 'neigh_op_lft_0')
// (8, 12, 'neigh_op_bnl_0')

wire n367;
// (6, 10, 'neigh_op_tnr_2')
// (6, 11, 'neigh_op_rgt_2')
// (6, 12, 'neigh_op_bnr_2')
// (7, 10, 'neigh_op_top_2')
// (7, 11, 'local_g2_2')
// (7, 11, 'lutff_1/in_3')
// (7, 11, 'lutff_2/out')
// (7, 12, 'neigh_op_bot_2')
// (8, 10, 'neigh_op_tnl_2')
// (8, 11, 'neigh_op_lft_2')
// (8, 12, 'neigh_op_bnl_2')

reg n368 = 0;
// (6, 10, 'neigh_op_tnr_3')
// (6, 11, 'neigh_op_rgt_3')
// (6, 12, 'neigh_op_bnr_3')
// (7, 10, 'neigh_op_top_3')
// (7, 11, 'local_g1_3')
// (7, 11, 'lutff_3/out')
// (7, 11, 'lutff_6/in_0')
// (7, 12, 'neigh_op_bot_3')
// (8, 10, 'neigh_op_tnl_3')
// (8, 11, 'neigh_op_lft_3')
// (8, 12, 'neigh_op_bnl_3')

reg n369 = 0;
// (6, 10, 'neigh_op_tnr_4')
// (6, 11, 'neigh_op_rgt_4')
// (6, 12, 'neigh_op_bnr_4')
// (7, 10, 'neigh_op_top_4')
// (7, 11, 'local_g0_4')
// (7, 11, 'lutff_0/in_2')
// (7, 11, 'lutff_4/out')
// (7, 11, 'lutff_7/in_1')
// (7, 12, 'neigh_op_bot_4')
// (8, 10, 'neigh_op_tnl_4')
// (8, 11, 'neigh_op_lft_4')
// (8, 12, 'neigh_op_bnl_4')

reg n370 = 0;
// (6, 10, 'neigh_op_tnr_5')
// (6, 11, 'neigh_op_rgt_5')
// (6, 12, 'neigh_op_bnr_5')
// (7, 10, 'neigh_op_top_5')
// (7, 11, 'local_g2_5')
// (7, 11, 'lutff_3/in_0')
// (7, 11, 'lutff_5/out')
// (7, 12, 'neigh_op_bot_5')
// (8, 10, 'neigh_op_tnl_5')
// (8, 11, 'neigh_op_lft_5')
// (8, 12, 'neigh_op_bnl_5')

reg n371 = 0;
// (6, 10, 'neigh_op_tnr_6')
// (6, 11, 'neigh_op_rgt_6')
// (6, 12, 'neigh_op_bnr_6')
// (7, 10, 'local_g1_6')
// (7, 10, 'lutff_3/in_0')
// (7, 10, 'neigh_op_top_6')
// (7, 11, 'lutff_6/out')
// (7, 12, 'local_g1_6')
// (7, 12, 'lutff_2/in_1')
// (7, 12, 'neigh_op_bot_6')
// (8, 10, 'neigh_op_tnl_6')
// (8, 11, 'neigh_op_lft_6')
// (8, 12, 'neigh_op_bnl_6')

wire n372;
// (6, 10, 'sp4_h_r_4')
// (6, 10, 'sp4_r_v_b_39')
// (6, 11, 'sp4_r_v_b_26')
// (6, 12, 'sp4_r_v_b_15')
// (6, 13, 'sp4_r_v_b_2')
// (7, 9, 'sp4_h_r_8')
// (7, 9, 'sp4_v_t_39')
// (7, 10, 'local_g0_1')
// (7, 10, 'lutff_0/in_1')
// (7, 10, 'sp4_h_r_17')
// (7, 10, 'sp4_v_b_39')
// (7, 11, 'sp4_v_b_26')
// (7, 12, 'sp4_v_b_15')
// (7, 13, 'local_g1_2')
// (7, 13, 'lutff_0/in_1')
// (7, 13, 'sp4_v_b_2')
// (8, 8, 'neigh_op_tnr_0')
// (8, 9, 'neigh_op_rgt_0')
// (8, 9, 'sp4_h_r_21')
// (8, 10, 'neigh_op_bnr_0')
// (8, 10, 'sp4_h_r_28')
// (9, 7, 'sp4_r_v_b_41')
// (9, 8, 'neigh_op_top_0')
// (9, 8, 'sp4_r_v_b_28')
// (9, 9, 'lutff_0/out')
// (9, 9, 'sp4_h_r_32')
// (9, 9, 'sp4_r_v_b_17')
// (9, 10, 'neigh_op_bot_0')
// (9, 10, 'sp4_h_r_41')
// (9, 10, 'sp4_r_v_b_4')
// (10, 6, 'sp4_v_t_41')
// (10, 7, 'sp4_v_b_41')
// (10, 8, 'neigh_op_tnl_0')
// (10, 8, 'sp4_v_b_28')
// (10, 9, 'neigh_op_lft_0')
// (10, 9, 'sp4_h_r_45')
// (10, 9, 'sp4_v_b_17')
// (10, 10, 'neigh_op_bnl_0')
// (10, 10, 'sp4_h_l_41')
// (10, 10, 'sp4_v_b_4')
// (11, 9, 'sp4_h_l_45')

reg n373 = 0;
// (6, 11, 'neigh_op_tnr_0')
// (6, 12, 'neigh_op_rgt_0')
// (6, 13, 'neigh_op_bnr_0')
// (7, 11, 'neigh_op_top_0')
// (7, 12, 'local_g0_0')
// (7, 12, 'lutff_0/out')
// (7, 12, 'lutff_6/in_0')
// (7, 13, 'neigh_op_bot_0')
// (8, 11, 'neigh_op_tnl_0')
// (8, 12, 'neigh_op_lft_0')
// (8, 13, 'neigh_op_bnl_0')

reg n374 = 0;
// (6, 11, 'neigh_op_tnr_1')
// (6, 12, 'neigh_op_rgt_1')
// (6, 13, 'neigh_op_bnr_1')
// (7, 11, 'neigh_op_top_1')
// (7, 12, 'local_g1_1')
// (7, 12, 'lutff_0/in_0')
// (7, 12, 'lutff_1/out')
// (7, 13, 'neigh_op_bot_1')
// (8, 11, 'neigh_op_tnl_1')
// (8, 12, 'neigh_op_lft_1')
// (8, 13, 'neigh_op_bnl_1')

reg n375 = 0;
// (6, 11, 'neigh_op_tnr_2')
// (6, 12, 'neigh_op_rgt_2')
// (6, 13, 'neigh_op_bnr_2')
// (7, 11, 'neigh_op_top_2')
// (7, 12, 'local_g1_2')
// (7, 12, 'lutff_1/in_0')
// (7, 12, 'lutff_2/out')
// (7, 13, 'neigh_op_bot_2')
// (8, 11, 'neigh_op_tnl_2')
// (8, 12, 'neigh_op_lft_2')
// (8, 13, 'neigh_op_bnl_2')

reg n376 = 0;
// (6, 11, 'neigh_op_tnr_3')
// (6, 12, 'neigh_op_rgt_3')
// (6, 13, 'neigh_op_bnr_3')
// (7, 11, 'neigh_op_top_3')
// (7, 12, 'lutff_3/out')
// (7, 13, 'local_g1_3')
// (7, 13, 'lutff_2/in_0')
// (7, 13, 'neigh_op_bot_3')
// (8, 11, 'neigh_op_tnl_3')
// (8, 12, 'neigh_op_lft_3')
// (8, 13, 'neigh_op_bnl_3')

reg n377 = 0;
// (6, 11, 'neigh_op_tnr_5')
// (6, 12, 'neigh_op_rgt_5')
// (6, 13, 'neigh_op_bnr_5')
// (7, 11, 'neigh_op_top_5')
// (7, 12, 'local_g0_5')
// (7, 12, 'lutff_5/out')
// (7, 12, 'lutff_7/in_0')
// (7, 13, 'neigh_op_bot_5')
// (8, 11, 'neigh_op_tnl_5')
// (8, 12, 'neigh_op_lft_5')
// (8, 13, 'neigh_op_bnl_5')

reg n378 = 0;
// (6, 11, 'neigh_op_tnr_7')
// (6, 12, 'neigh_op_rgt_7')
// (6, 13, 'neigh_op_bnr_7')
// (7, 11, 'neigh_op_top_7')
// (7, 12, 'lutff_7/out')
// (7, 13, 'neigh_op_bot_7')
// (8, 11, 'neigh_op_tnl_7')
// (8, 12, 'local_g1_7')
// (8, 12, 'lutff_6/in_0')
// (8, 12, 'neigh_op_lft_7')
// (8, 13, 'neigh_op_bnl_7')

reg n379 = 0;
// (6, 11, 'sp4_h_r_0')
// (7, 10, 'neigh_op_tnr_4')
// (7, 11, 'local_g0_5')
// (7, 11, 'lutff_0/in_1')
// (7, 11, 'neigh_op_rgt_4')
// (7, 11, 'sp4_h_r_13')
// (7, 12, 'neigh_op_bnr_4')
// (8, 10, 'neigh_op_top_4')
// (8, 11, 'lutff_4/out')
// (8, 11, 'sp4_h_r_24')
// (8, 12, 'neigh_op_bot_4')
// (9, 10, 'neigh_op_tnl_4')
// (9, 11, 'neigh_op_lft_4')
// (9, 11, 'sp4_h_r_37')
// (9, 12, 'neigh_op_bnl_4')
// (10, 11, 'sp4_h_l_37')

reg n380 = 0;
// (6, 11, 'sp4_r_v_b_36')
// (6, 12, 'local_g1_1')
// (6, 12, 'lutff_2/in_0')
// (6, 12, 'neigh_op_tnr_6')
// (6, 12, 'sp4_r_v_b_25')
// (6, 13, 'neigh_op_rgt_6')
// (6, 13, 'sp4_r_v_b_12')
// (6, 14, 'neigh_op_bnr_6')
// (6, 14, 'sp4_r_v_b_1')
// (7, 10, 'sp4_v_t_36')
// (7, 11, 'sp4_v_b_36')
// (7, 12, 'neigh_op_top_6')
// (7, 12, 'sp4_v_b_25')
// (7, 13, 'local_g0_6')
// (7, 13, 'lutff_3/in_1')
// (7, 13, 'lutff_6/out')
// (7, 13, 'sp4_v_b_12')
// (7, 14, 'neigh_op_bot_6')
// (7, 14, 'sp4_v_b_1')
// (8, 12, 'neigh_op_tnl_6')
// (8, 13, 'neigh_op_lft_6')
// (8, 14, 'neigh_op_bnl_6')

reg n381 = 0;
// (6, 12, 'neigh_op_tnr_0')
// (6, 13, 'neigh_op_rgt_0')
// (6, 14, 'neigh_op_bnr_0')
// (7, 12, 'neigh_op_top_0')
// (7, 13, 'local_g1_0')
// (7, 13, 'lutff_0/out')
// (7, 13, 'lutff_5/in_0')
// (7, 14, 'neigh_op_bot_0')
// (8, 12, 'neigh_op_tnl_0')
// (8, 13, 'neigh_op_lft_0')
// (8, 14, 'neigh_op_bnl_0')

reg n382 = 0;
// (6, 12, 'neigh_op_tnr_2')
// (6, 13, 'neigh_op_rgt_2')
// (6, 14, 'neigh_op_bnr_2')
// (7, 12, 'neigh_op_top_2')
// (7, 13, 'local_g0_2')
// (7, 13, 'lutff_2/out')
// (7, 13, 'lutff_6/in_0')
// (7, 14, 'neigh_op_bot_2')
// (8, 12, 'neigh_op_tnl_2')
// (8, 13, 'neigh_op_lft_2')
// (8, 14, 'neigh_op_bnl_2')

reg n383 = 0;
// (6, 12, 'neigh_op_tnr_3')
// (6, 13, 'neigh_op_rgt_3')
// (6, 14, 'neigh_op_bnr_3')
// (7, 12, 'neigh_op_top_3')
// (7, 13, 'lutff_3/out')
// (7, 13, 'sp4_h_r_6')
// (7, 14, 'neigh_op_bot_3')
// (8, 12, 'neigh_op_tnl_3')
// (8, 13, 'neigh_op_lft_3')
// (8, 13, 'sp4_h_r_19')
// (8, 14, 'neigh_op_bnl_3')
// (9, 13, 'sp4_h_r_30')
// (10, 13, 'sp4_h_r_43')
// (11, 13, 'local_g0_1')
// (11, 13, 'lutff_7/in_0')
// (11, 13, 'sp4_h_l_43')
// (11, 13, 'sp4_h_r_9')
// (12, 13, 'sp4_h_r_20')
// (13, 13, 'span4_horz_20')

reg n384 = 0;
// (6, 12, 'neigh_op_tnr_4')
// (6, 13, 'neigh_op_rgt_4')
// (6, 14, 'neigh_op_bnr_4')
// (7, 12, 'neigh_op_top_4')
// (7, 13, 'local_g1_4')
// (7, 13, 'lutff_4/out')
// (7, 13, 'lutff_7/in_0')
// (7, 14, 'neigh_op_bot_4')
// (8, 12, 'neigh_op_tnl_4')
// (8, 13, 'neigh_op_lft_4')
// (8, 14, 'neigh_op_bnl_4')

reg n385 = 0;
// (6, 12, 'neigh_op_tnr_5')
// (6, 13, 'neigh_op_rgt_5')
// (6, 14, 'neigh_op_bnr_5')
// (7, 12, 'neigh_op_top_5')
// (7, 13, 'local_g1_5')
// (7, 13, 'lutff_4/in_0')
// (7, 13, 'lutff_5/out')
// (7, 14, 'neigh_op_bot_5')
// (8, 12, 'neigh_op_tnl_5')
// (8, 13, 'neigh_op_lft_5')
// (8, 14, 'neigh_op_bnl_5')

reg n386 = 0;
// (6, 12, 'neigh_op_tnr_7')
// (6, 13, 'neigh_op_rgt_7')
// (6, 14, 'neigh_op_bnr_7')
// (7, 12, 'neigh_op_top_7')
// (7, 13, 'lutff_7/out')
// (7, 14, 'local_g0_7')
// (7, 14, 'local_g1_7')
// (7, 14, 'lutff_0/in_1')
// (7, 14, 'lutff_5/in_1')
// (7, 14, 'neigh_op_bot_7')
// (8, 12, 'neigh_op_tnl_7')
// (8, 13, 'neigh_op_lft_7')
// (8, 14, 'neigh_op_bnl_7')

reg n387 = 0;
// (6, 12, 'sp12_h_r_1')
// (7, 12, 'sp12_h_r_2')
// (8, 12, 'local_g0_5')
// (8, 12, 'lutff_1/in_2')
// (8, 12, 'sp12_h_r_5')
// (9, 12, 'local_g1_6')
// (9, 12, 'lutff_6/in_1')
// (9, 12, 'sp12_h_r_6')
// (10, 11, 'neigh_op_tnr_1')
// (10, 12, 'neigh_op_rgt_1')
// (10, 12, 'sp12_h_r_9')
// (10, 13, 'neigh_op_bnr_1')
// (11, 11, 'neigh_op_top_1')
// (11, 12, 'lutff_1/out')
// (11, 12, 'sp12_h_r_10')
// (11, 13, 'neigh_op_bot_1')
// (12, 11, 'neigh_op_tnl_1')
// (12, 12, 'neigh_op_lft_1')
// (12, 12, 'sp12_h_r_13')
// (12, 13, 'neigh_op_bnl_1')
// (13, 12, 'span12_horz_13')

wire n388;
// (6, 13, 'neigh_op_tnr_0')
// (6, 14, 'neigh_op_rgt_0')
// (6, 15, 'neigh_op_bnr_0')
// (7, 13, 'neigh_op_top_0')
// (7, 13, 'sp4_r_v_b_44')
// (7, 14, 'local_g0_2')
// (7, 14, 'lutff_0/out')
// (7, 14, 'lutff_1/in_3')
// (7, 14, 'sp4_r_v_b_33')
// (7, 15, 'neigh_op_bot_0')
// (7, 15, 'sp4_r_v_b_20')
// (7, 16, 'sp4_r_v_b_9')
// (8, 12, 'sp4_v_t_44')
// (8, 13, 'neigh_op_tnl_0')
// (8, 13, 'sp4_v_b_44')
// (8, 14, 'neigh_op_lft_0')
// (8, 14, 'sp4_v_b_33')
// (8, 15, 'neigh_op_bnl_0')
// (8, 15, 'sp4_v_b_20')
// (8, 16, 'sp4_v_b_9')

wire n389;
// (6, 13, 'neigh_op_tnr_1')
// (6, 14, 'neigh_op_rgt_1')
// (6, 15, 'neigh_op_bnr_1')
// (7, 3, 'sp12_v_t_22')
// (7, 4, 'sp12_v_b_22')
// (7, 5, 'sp12_v_b_21')
// (7, 6, 'sp12_v_b_18')
// (7, 7, 'sp12_v_b_17')
// (7, 8, 'sp12_v_b_14')
// (7, 9, 'sp12_v_b_13')
// (7, 10, 'local_g3_2')
// (7, 10, 'lutff_0/in_3')
// (7, 10, 'sp12_v_b_10')
// (7, 11, 'sp12_v_b_9')
// (7, 12, 'sp12_v_b_6')
// (7, 13, 'neigh_op_top_1')
// (7, 13, 'sp12_v_b_5')
// (7, 14, 'lutff_1/out')
// (7, 14, 'sp12_v_b_2')
// (7, 15, 'neigh_op_bot_1')
// (7, 15, 'sp12_v_b_1')
// (8, 13, 'neigh_op_tnl_1')
// (8, 14, 'neigh_op_lft_1')
// (8, 15, 'neigh_op_bnl_1')

reg n390 = 0;
// (6, 13, 'neigh_op_tnr_2')
// (6, 14, 'neigh_op_rgt_2')
// (6, 15, 'neigh_op_bnr_2')
// (7, 13, 'neigh_op_top_2')
// (7, 14, 'lutff_2/out')
// (7, 15, 'local_g1_2')
// (7, 15, 'lutff_7/in_0')
// (7, 15, 'neigh_op_bot_2')
// (8, 13, 'neigh_op_tnl_2')
// (8, 14, 'neigh_op_lft_2')
// (8, 15, 'neigh_op_bnl_2')

reg n391 = 0;
// (6, 13, 'neigh_op_tnr_3')
// (6, 14, 'neigh_op_rgt_3')
// (6, 15, 'neigh_op_bnr_3')
// (7, 13, 'neigh_op_top_3')
// (7, 14, 'local_g1_3')
// (7, 14, 'lutff_3/out')
// (7, 14, 'lutff_4/in_0')
// (7, 15, 'neigh_op_bot_3')
// (8, 13, 'neigh_op_tnl_3')
// (8, 14, 'neigh_op_lft_3')
// (8, 15, 'neigh_op_bnl_3')

reg n392 = 0;
// (6, 13, 'neigh_op_tnr_4')
// (6, 14, 'neigh_op_rgt_4')
// (6, 15, 'neigh_op_bnr_4')
// (7, 13, 'neigh_op_top_4')
// (7, 14, 'local_g0_4')
// (7, 14, 'local_g1_4')
// (7, 14, 'lutff_0/in_0')
// (7, 14, 'lutff_2/in_1')
// (7, 14, 'lutff_4/out')
// (7, 15, 'neigh_op_bot_4')
// (8, 13, 'neigh_op_tnl_4')
// (8, 14, 'neigh_op_lft_4')
// (8, 15, 'neigh_op_bnl_4')

reg n393 = 0;
// (6, 13, 'neigh_op_tnr_5')
// (6, 14, 'neigh_op_rgt_5')
// (6, 15, 'neigh_op_bnr_5')
// (7, 13, 'neigh_op_top_5')
// (7, 14, 'local_g1_5')
// (7, 14, 'lutff_5/out')
// (7, 14, 'lutff_6/in_0')
// (7, 15, 'neigh_op_bot_5')
// (8, 13, 'neigh_op_tnl_5')
// (8, 14, 'neigh_op_lft_5')
// (8, 15, 'neigh_op_bnl_5')

reg n394 = 0;
// (6, 13, 'neigh_op_tnr_6')
// (6, 14, 'neigh_op_rgt_6')
// (6, 15, 'neigh_op_bnr_6')
// (7, 13, 'neigh_op_top_6')
// (7, 14, 'local_g1_6')
// (7, 14, 'lutff_3/in_0')
// (7, 14, 'lutff_6/out')
// (7, 15, 'neigh_op_bot_6')
// (8, 13, 'neigh_op_tnl_6')
// (8, 14, 'neigh_op_lft_6')
// (8, 15, 'neigh_op_bnl_6')

reg n395 = 0;
// (6, 14, 'neigh_op_tnr_2')
// (6, 15, 'neigh_op_rgt_2')
// (6, 16, 'neigh_op_bnr_2')
// (7, 5, 'sp12_v_t_23')
// (7, 6, 'sp12_v_b_23')
// (7, 7, 'sp12_v_b_20')
// (7, 8, 'sp12_v_b_19')
// (7, 9, 'sp12_v_b_16')
// (7, 10, 'sp12_v_b_15')
// (7, 11, 'sp12_v_b_12')
// (7, 12, 'sp12_v_b_11')
// (7, 13, 'local_g2_0')
// (7, 13, 'lutff_0/in_0')
// (7, 13, 'sp12_v_b_8')
// (7, 14, 'local_g1_2')
// (7, 14, 'local_g3_7')
// (7, 14, 'lutff_1/in_0')
// (7, 14, 'lutff_2/in_0')
// (7, 14, 'lutff_5/in_0')
// (7, 14, 'neigh_op_top_2')
// (7, 14, 'sp12_v_b_7')
// (7, 15, 'lutff_2/out')
// (7, 15, 'sp12_v_b_4')
// (7, 16, 'neigh_op_bot_2')
// (7, 16, 'sp12_v_b_3')
// (7, 17, 'span12_vert_0')
// (8, 14, 'neigh_op_tnl_2')
// (8, 15, 'neigh_op_lft_2')
// (8, 16, 'neigh_op_bnl_2')

reg n396 = 0;
// (6, 14, 'neigh_op_tnr_4')
// (6, 15, 'neigh_op_rgt_4')
// (6, 16, 'neigh_op_bnr_4')
// (7, 14, 'neigh_op_top_4')
// (7, 15, 'local_g0_4')
// (7, 15, 'lutff_2/in_0')
// (7, 15, 'lutff_4/out')
// (7, 16, 'neigh_op_bot_4')
// (8, 14, 'neigh_op_tnl_4')
// (8, 15, 'neigh_op_lft_4')
// (8, 16, 'neigh_op_bnl_4')

reg n397 = 0;
// (6, 14, 'neigh_op_tnr_7')
// (6, 15, 'neigh_op_rgt_7')
// (6, 16, 'neigh_op_bnr_7')
// (7, 14, 'neigh_op_top_7')
// (7, 15, 'local_g1_7')
// (7, 15, 'lutff_4/in_0')
// (7, 15, 'lutff_7/out')
// (7, 16, 'neigh_op_bot_7')
// (8, 14, 'neigh_op_tnl_7')
// (8, 15, 'neigh_op_lft_7')
// (8, 16, 'neigh_op_bnl_7')

wire n398;
// (7, 1, 'neigh_op_tnr_0')
// (7, 2, 'neigh_op_rgt_0')
// (7, 3, 'neigh_op_bnr_0')
// (8, 1, 'neigh_op_top_0')
// (8, 2, 'local_g1_0')
// (8, 2, 'local_g2_0')
// (8, 2, 'lutff_0/out')
// (8, 2, 'lutff_1/in_3')
// (8, 2, 'lutff_2/in_1')
// (8, 2, 'lutff_3/in_1')
// (8, 2, 'lutff_4/in_0')
// (8, 2, 'lutff_5/in_3')
// (8, 2, 'lutff_6/in_3')
// (8, 2, 'lutff_7/in_3')
// (8, 3, 'neigh_op_bot_0')
// (9, 1, 'neigh_op_tnl_0')
// (9, 2, 'neigh_op_lft_0')
// (9, 3, 'neigh_op_bnl_0')

wire n399;
// (7, 1, 'neigh_op_tnr_1')
// (7, 1, 'sp4_r_v_b_47')
// (7, 2, 'neigh_op_rgt_1')
// (7, 2, 'sp4_r_v_b_34')
// (7, 3, 'neigh_op_bnr_1')
// (7, 3, 'sp4_r_v_b_23')
// (7, 4, 'sp4_r_v_b_10')
// (8, 0, 'span4_vert_47')
// (8, 1, 'neigh_op_top_1')
// (8, 1, 'sp4_v_b_47')
// (8, 2, 'lutff_1/out')
// (8, 2, 'sp4_v_b_34')
// (8, 3, 'local_g0_1')
// (8, 3, 'lutff_6/in_1')
// (8, 3, 'neigh_op_bot_1')
// (8, 3, 'sp4_v_b_23')
// (8, 4, 'local_g1_2')
// (8, 4, 'lutff_2/in_1')
// (8, 4, 'sp4_v_b_10')
// (9, 1, 'neigh_op_tnl_1')
// (9, 2, 'neigh_op_lft_1')
// (9, 3, 'neigh_op_bnl_1')

wire n400;
// (7, 1, 'neigh_op_tnr_2')
// (7, 2, 'neigh_op_rgt_2')
// (7, 3, 'neigh_op_bnr_2')
// (8, 1, 'neigh_op_top_2')
// (8, 2, 'lutff_2/out')
// (8, 3, 'local_g1_2')
// (8, 3, 'lutff_3/in_0')
// (8, 3, 'lutff_5/in_0')
// (8, 3, 'neigh_op_bot_2')
// (9, 1, 'neigh_op_tnl_2')
// (9, 2, 'neigh_op_lft_2')
// (9, 3, 'neigh_op_bnl_2')

wire n401;
// (7, 1, 'neigh_op_tnr_3')
// (7, 2, 'neigh_op_rgt_3')
// (7, 3, 'neigh_op_bnr_3')
// (7, 3, 'sp4_r_v_b_36')
// (7, 4, 'local_g0_1')
// (7, 4, 'lutff_1/in_0')
// (7, 4, 'sp4_r_v_b_25')
// (7, 5, 'sp4_r_v_b_12')
// (7, 6, 'sp4_r_v_b_1')
// (8, 0, 'span12_vert_9')
// (8, 1, 'neigh_op_top_3')
// (8, 1, 'sp12_v_b_9')
// (8, 2, 'lutff_3/out')
// (8, 2, 'sp12_v_b_6')
// (8, 2, 'sp4_v_t_36')
// (8, 3, 'local_g0_3')
// (8, 3, 'lutff_4/in_1')
// (8, 3, 'neigh_op_bot_3')
// (8, 3, 'sp12_v_b_5')
// (8, 3, 'sp4_v_b_36')
// (8, 4, 'sp12_v_b_2')
// (8, 4, 'sp4_v_b_25')
// (8, 5, 'sp12_v_b_1')
// (8, 5, 'sp4_v_b_12')
// (8, 6, 'sp4_v_b_1')
// (9, 1, 'neigh_op_tnl_3')
// (9, 2, 'neigh_op_lft_3')
// (9, 3, 'neigh_op_bnl_3')

wire n402;
// (7, 1, 'neigh_op_tnr_4')
// (7, 2, 'neigh_op_rgt_4')
// (7, 3, 'neigh_op_bnr_4')
// (8, 1, 'neigh_op_top_4')
// (8, 2, 'lutff_4/out')
// (8, 3, 'local_g0_4')
// (8, 3, 'lutff_0/in_0')
// (8, 3, 'lutff_2/in_0')
// (8, 3, 'neigh_op_bot_4')
// (9, 1, 'neigh_op_tnl_4')
// (9, 2, 'neigh_op_lft_4')
// (9, 3, 'neigh_op_bnl_4')

wire n403;
// (7, 1, 'neigh_op_tnr_6')
// (7, 1, 'sp4_r_v_b_41')
// (7, 2, 'neigh_op_rgt_6')
// (7, 2, 'sp4_r_v_b_28')
// (7, 3, 'neigh_op_bnr_6')
// (7, 3, 'sp4_r_v_b_17')
// (7, 4, 'sp4_r_v_b_4')
// (8, 0, 'span4_vert_41')
// (8, 1, 'neigh_op_top_6')
// (8, 1, 'sp4_v_b_41')
// (8, 2, 'lutff_6/out')
// (8, 2, 'sp4_v_b_28')
// (8, 3, 'local_g0_6')
// (8, 3, 'lutff_7/in_1')
// (8, 3, 'neigh_op_bot_6')
// (8, 3, 'sp4_v_b_17')
// (8, 4, 'local_g0_4')
// (8, 4, 'local_g1_4')
// (8, 4, 'lutff_4/in_1')
// (8, 4, 'lutff_5/in_2')
// (8, 4, 'lutff_7/in_1')
// (8, 4, 'sp4_v_b_4')
// (9, 1, 'neigh_op_tnl_6')
// (9, 2, 'neigh_op_lft_6')
// (9, 3, 'neigh_op_bnl_6')

wire n404;
// (7, 1, 'neigh_op_tnr_7')
// (7, 2, 'neigh_op_rgt_7')
// (7, 3, 'neigh_op_bnr_7')
// (8, 1, 'neigh_op_top_7')
// (8, 2, 'lutff_7/out')
// (8, 3, 'local_g0_7')
// (8, 3, 'local_g1_7')
// (8, 3, 'lutff_0/in_2')
// (8, 3, 'lutff_2/in_2')
// (8, 3, 'lutff_3/in_2')
// (8, 3, 'lutff_5/in_2')
// (8, 3, 'neigh_op_bot_7')
// (9, 1, 'neigh_op_tnl_7')
// (9, 2, 'neigh_op_lft_7')
// (9, 3, 'neigh_op_bnl_7')

wire n405;
// (7, 1, 'sp4_r_v_b_44')
// (7, 2, 'neigh_op_tnr_2')
// (7, 2, 'sp4_r_v_b_33')
// (7, 3, 'neigh_op_rgt_2')
// (7, 3, 'sp4_r_v_b_20')
// (7, 4, 'neigh_op_bnr_2')
// (7, 4, 'sp4_r_v_b_9')
// (8, 0, 'span4_vert_44')
// (8, 1, 'sp4_v_b_44')
// (8, 2, 'neigh_op_top_2')
// (8, 2, 'sp4_v_b_33')
// (8, 3, 'lutff_2/out')
// (8, 3, 'sp4_v_b_20')
// (8, 4, 'local_g1_1')
// (8, 4, 'lutff_1/in_3')
// (8, 4, 'neigh_op_bot_2')
// (8, 4, 'sp4_v_b_9')
// (9, 2, 'neigh_op_tnl_2')
// (9, 3, 'neigh_op_lft_2')
// (9, 4, 'neigh_op_bnl_2')

wire n406;
// (7, 2, 'local_g3_1')
// (7, 2, 'lutff_2/in_2')
// (7, 2, 'lutff_5/in_1')
// (7, 2, 'neigh_op_tnr_1')
// (7, 3, 'neigh_op_rgt_1')
// (7, 4, 'neigh_op_bnr_1')
// (8, 2, 'local_g1_1')
// (8, 2, 'lutff_0/in_2')
// (8, 2, 'neigh_op_top_1')
// (8, 3, 'lutff_1/out')
// (8, 4, 'neigh_op_bot_1')
// (9, 2, 'neigh_op_tnl_1')
// (9, 3, 'neigh_op_lft_1')
// (9, 4, 'neigh_op_bnl_1')

wire n407;
// (7, 2, 'neigh_op_tnr_3')
// (7, 3, 'neigh_op_rgt_3')
// (7, 4, 'neigh_op_bnr_3')
// (8, 0, 'span12_vert_10')
// (8, 1, 'sp12_v_b_10')
// (8, 2, 'neigh_op_top_3')
// (8, 2, 'sp12_v_b_9')
// (8, 3, 'lutff_3/out')
// (8, 3, 'sp12_v_b_6')
// (8, 4, 'neigh_op_bot_3')
// (8, 4, 'sp12_v_b_5')
// (8, 5, 'local_g2_2')
// (8, 5, 'lutff_7/in_3')
// (8, 5, 'sp12_v_b_2')
// (8, 6, 'sp12_v_b_1')
// (9, 2, 'neigh_op_tnl_3')
// (9, 3, 'neigh_op_lft_3')
// (9, 4, 'neigh_op_bnl_3')

wire n408;
// (7, 2, 'neigh_op_tnr_4')
// (7, 3, 'neigh_op_rgt_4')
// (7, 4, 'neigh_op_bnr_4')
// (7, 4, 'sp4_r_v_b_37')
// (7, 5, 'sp4_r_v_b_24')
// (7, 6, 'sp4_r_v_b_13')
// (7, 7, 'sp4_r_v_b_0')
// (8, 0, 'span12_vert_12')
// (8, 1, 'sp12_v_b_12')
// (8, 2, 'neigh_op_top_4')
// (8, 2, 'sp12_v_b_11')
// (8, 3, 'lutff_4/out')
// (8, 3, 'sp12_v_b_8')
// (8, 3, 'sp4_v_t_37')
// (8, 4, 'local_g2_7')
// (8, 4, 'lutff_1/in_0')
// (8, 4, 'neigh_op_bot_4')
// (8, 4, 'sp12_v_b_7')
// (8, 4, 'sp4_v_b_37')
// (8, 5, 'local_g2_0')
// (8, 5, 'lutff_2/in_2')
// (8, 5, 'lutff_5/in_1')
// (8, 5, 'sp12_v_b_4')
// (8, 5, 'sp4_v_b_24')
// (8, 6, 'sp12_v_b_3')
// (8, 6, 'sp4_v_b_13')
// (8, 7, 'sp12_v_b_0')
// (8, 7, 'sp4_v_b_0')
// (9, 2, 'neigh_op_tnl_4')
// (9, 3, 'neigh_op_lft_4')
// (9, 4, 'neigh_op_bnl_4')

wire n409;
// (7, 2, 'neigh_op_tnr_5')
// (7, 3, 'neigh_op_rgt_5')
// (7, 4, 'neigh_op_bnr_5')
// (8, 2, 'neigh_op_top_5')
// (8, 2, 'sp4_r_v_b_38')
// (8, 3, 'lutff_5/out')
// (8, 3, 'sp4_r_v_b_27')
// (8, 3, 'sp4_r_v_b_43')
// (8, 4, 'local_g1_6')
// (8, 4, 'local_g2_6')
// (8, 4, 'lutff_0/in_3')
// (8, 4, 'lutff_6/in_2')
// (8, 4, 'neigh_op_bot_5')
// (8, 4, 'sp4_r_v_b_14')
// (8, 4, 'sp4_r_v_b_30')
// (8, 5, 'sp4_r_v_b_19')
// (8, 5, 'sp4_r_v_b_3')
// (8, 6, 'sp4_r_v_b_6')
// (9, 1, 'sp4_v_t_38')
// (9, 2, 'neigh_op_tnl_5')
// (9, 2, 'sp4_v_b_38')
// (9, 2, 'sp4_v_t_43')
// (9, 3, 'neigh_op_lft_5')
// (9, 3, 'sp4_v_b_27')
// (9, 3, 'sp4_v_b_43')
// (9, 4, 'neigh_op_bnl_5')
// (9, 4, 'sp4_v_b_14')
// (9, 4, 'sp4_v_b_30')
// (9, 5, 'sp4_v_b_19')
// (9, 5, 'sp4_v_b_3')
// (9, 6, 'sp4_v_b_6')

wire n410;
// (7, 2, 'neigh_op_tnr_7')
// (7, 3, 'neigh_op_rgt_7')
// (7, 4, 'neigh_op_bnr_7')
// (8, 2, 'neigh_op_top_7')
// (8, 3, 'local_g3_7')
// (8, 3, 'lutff_6/in_2')
// (8, 3, 'lutff_7/out')
// (8, 3, 'sp4_r_v_b_47')
// (8, 4, 'local_g0_1')
// (8, 4, 'local_g1_7')
// (8, 4, 'lutff_0/in_2')
// (8, 4, 'lutff_6/in_1')
// (8, 4, 'neigh_op_bot_7')
// (8, 4, 'sp4_r_v_b_34')
// (8, 5, 'sp4_r_v_b_23')
// (8, 6, 'sp4_r_v_b_10')
// (9, 2, 'neigh_op_tnl_7')
// (9, 2, 'sp4_v_t_47')
// (9, 3, 'neigh_op_lft_7')
// (9, 3, 'sp4_v_b_47')
// (9, 4, 'neigh_op_bnl_7')
// (9, 4, 'sp4_v_b_34')
// (9, 5, 'sp4_v_b_23')
// (9, 6, 'sp4_v_b_10')

wire n411;
// (7, 2, 'sp4_r_v_b_38')
// (7, 3, 'neigh_op_tnr_7')
// (7, 3, 'sp4_r_v_b_27')
// (7, 4, 'neigh_op_rgt_7')
// (7, 4, 'sp4_r_v_b_14')
// (7, 5, 'neigh_op_bnr_7')
// (7, 5, 'sp4_r_v_b_3')
// (8, 1, 'sp4_v_t_38')
// (8, 2, 'sp4_v_b_38')
// (8, 3, 'neigh_op_top_7')
// (8, 3, 'sp4_v_b_27')
// (8, 4, 'local_g3_7')
// (8, 4, 'lutff_1/in_1')
// (8, 4, 'lutff_7/out')
// (8, 4, 'sp4_v_b_14')
// (8, 5, 'local_g0_3')
// (8, 5, 'lutff_6/in_3')
// (8, 5, 'neigh_op_bot_7')
// (8, 5, 'sp4_v_b_3')
// (9, 3, 'neigh_op_tnl_7')
// (9, 4, 'neigh_op_lft_7')
// (9, 5, 'neigh_op_bnl_7')

wire n412;
// (7, 3, 'neigh_op_tnr_0')
// (7, 4, 'neigh_op_rgt_0')
// (7, 5, 'neigh_op_bnr_0')
// (8, 3, 'neigh_op_top_0')
// (8, 4, 'lutff_0/out')
// (8, 5, 'local_g1_0')
// (8, 5, 'lutff_0/in_1')
// (8, 5, 'neigh_op_bot_0')
// (9, 3, 'neigh_op_tnl_0')
// (9, 4, 'neigh_op_lft_0')
// (9, 5, 'neigh_op_bnl_0')

wire n413;
// (7, 3, 'neigh_op_tnr_1')
// (7, 3, 'sp4_r_v_b_47')
// (7, 4, 'neigh_op_rgt_1')
// (7, 4, 'sp4_r_v_b_34')
// (7, 5, 'local_g0_1')
// (7, 5, 'lutff_6/in_1')
// (7, 5, 'neigh_op_bnr_1')
// (7, 5, 'sp4_r_v_b_23')
// (7, 6, 'local_g2_2')
// (7, 6, 'lutff_5/in_1')
// (7, 6, 'sp4_r_v_b_10')
// (8, 2, 'sp4_v_t_47')
// (8, 3, 'neigh_op_top_1')
// (8, 3, 'sp4_v_b_47')
// (8, 4, 'lutff_1/out')
// (8, 4, 'sp4_v_b_34')
// (8, 5, 'neigh_op_bot_1')
// (8, 5, 'sp4_v_b_23')
// (8, 6, 'sp4_v_b_10')
// (9, 3, 'neigh_op_tnl_1')
// (9, 4, 'neigh_op_lft_1')
// (9, 5, 'neigh_op_bnl_1')

wire n414;
// (7, 3, 'neigh_op_tnr_2')
// (7, 4, 'neigh_op_rgt_2')
// (7, 5, 'neigh_op_bnr_2')
// (8, 3, 'neigh_op_top_2')
// (8, 4, 'local_g0_2')
// (8, 4, 'local_g3_2')
// (8, 4, 'lutff_2/out')
// (8, 4, 'lutff_3/in_3')
// (8, 4, 'lutff_6/in_3')
// (8, 5, 'neigh_op_bot_2')
// (9, 3, 'neigh_op_tnl_2')
// (9, 4, 'neigh_op_lft_2')
// (9, 5, 'neigh_op_bnl_2')

wire n415;
// (7, 3, 'neigh_op_tnr_4')
// (7, 4, 'local_g3_4')
// (7, 4, 'lutff_1/in_2')
// (7, 4, 'neigh_op_rgt_4')
// (7, 5, 'neigh_op_bnr_4')
// (8, 3, 'neigh_op_top_4')
// (8, 4, 'local_g3_4')
// (8, 4, 'lutff_1/in_2')
// (8, 4, 'lutff_4/out')
// (8, 5, 'neigh_op_bot_4')
// (9, 3, 'neigh_op_tnl_4')
// (9, 4, 'neigh_op_lft_4')
// (9, 5, 'neigh_op_bnl_4')

wire n416;
// (7, 3, 'neigh_op_tnr_5')
// (7, 4, 'neigh_op_rgt_5')
// (7, 5, 'neigh_op_bnr_5')
// (8, 3, 'neigh_op_top_5')
// (8, 4, 'local_g0_5')
// (8, 4, 'local_g1_5')
// (8, 4, 'lutff_3/in_2')
// (8, 4, 'lutff_5/out')
// (8, 4, 'lutff_6/in_0')
// (8, 4, 'sp4_r_v_b_43')
// (8, 5, 'local_g1_6')
// (8, 5, 'lutff_7/in_2')
// (8, 5, 'neigh_op_bot_5')
// (8, 5, 'sp4_r_v_b_30')
// (8, 6, 'sp4_r_v_b_19')
// (8, 7, 'sp4_r_v_b_6')
// (9, 3, 'neigh_op_tnl_5')
// (9, 3, 'sp4_v_t_43')
// (9, 4, 'neigh_op_lft_5')
// (9, 4, 'sp4_v_b_43')
// (9, 5, 'neigh_op_bnl_5')
// (9, 5, 'sp4_v_b_30')
// (9, 6, 'sp4_v_b_19')
// (9, 7, 'sp4_v_b_6')

reg n417 = 0;
// (7, 3, 'sp4_r_v_b_37')
// (7, 4, 'sp4_r_v_b_24')
// (7, 5, 'local_g2_5')
// (7, 5, 'lutff_1/in_2')
// (7, 5, 'sp4_r_v_b_13')
// (7, 6, 'sp4_r_v_b_0')
// (8, 2, 'sp4_v_t_37')
// (8, 3, 'sp4_v_b_37')
// (8, 4, 'sp4_v_b_24')
// (8, 5, 'sp4_v_b_13')
// (8, 6, 'sp4_h_r_7')
// (8, 6, 'sp4_v_b_0')
// (9, 6, 'sp4_h_r_18')
// (10, 5, 'neigh_op_tnr_5')
// (10, 6, 'neigh_op_rgt_5')
// (10, 6, 'sp4_h_r_31')
// (10, 7, 'neigh_op_bnr_5')
// (11, 5, 'neigh_op_top_5')
// (11, 6, 'local_g1_5')
// (11, 6, 'lutff_4/in_0')
// (11, 6, 'lutff_5/out')
// (11, 6, 'sp4_h_r_42')
// (11, 7, 'neigh_op_bot_5')
// (12, 5, 'neigh_op_tnl_5')
// (12, 6, 'neigh_op_lft_5')
// (12, 6, 'sp4_h_l_42')
// (12, 7, 'neigh_op_bnl_5')

wire n418;
// (7, 4, 'neigh_op_tnr_0')
// (7, 5, 'neigh_op_rgt_0')
// (7, 6, 'neigh_op_bnr_0')
// (8, 2, 'sp4_r_v_b_36')
// (8, 3, 'sp4_r_v_b_25')
// (8, 4, 'neigh_op_top_0')
// (8, 4, 'sp4_r_v_b_12')
// (8, 5, 'lutff_0/out')
// (8, 5, 'sp4_r_v_b_1')
// (8, 6, 'neigh_op_bot_0')
// (8, 6, 'sp4_r_v_b_36')
// (8, 7, 'sp4_r_v_b_25')
// (8, 8, 'sp4_r_v_b_12')
// (8, 9, 'sp4_r_v_b_1')
// (9, 1, 'sp4_v_t_36')
// (9, 2, 'sp4_v_b_36')
// (9, 3, 'sp4_v_b_25')
// (9, 4, 'neigh_op_tnl_0')
// (9, 4, 'sp4_v_b_12')
// (9, 5, 'neigh_op_lft_0')
// (9, 5, 'sp4_v_b_1')
// (9, 5, 'sp4_v_t_36')
// (9, 6, 'local_g2_0')
// (9, 6, 'lutff_6/in_2')
// (9, 6, 'neigh_op_bnl_0')
// (9, 6, 'sp4_v_b_36')
// (9, 7, 'sp4_v_b_25')
// (9, 8, 'local_g0_4')
// (9, 8, 'lutff_3/in_1')
// (9, 8, 'lutff_5/in_1')
// (9, 8, 'sp4_v_b_12')
// (9, 9, 'sp4_v_b_1')

wire n419;
// (7, 4, 'neigh_op_tnr_2')
// (7, 5, 'neigh_op_rgt_2')
// (7, 6, 'neigh_op_bnr_2')
// (8, 4, 'neigh_op_top_2')
// (8, 5, 'local_g1_2')
// (8, 5, 'lutff_2/out')
// (8, 5, 'lutff_4/in_1')
// (8, 6, 'neigh_op_bot_2')
// (9, 4, 'neigh_op_tnl_2')
// (9, 5, 'neigh_op_lft_2')
// (9, 6, 'neigh_op_bnl_2')

wire n420;
// (7, 4, 'neigh_op_tnr_3')
// (7, 5, 'neigh_op_rgt_3')
// (7, 6, 'neigh_op_bnr_3')
// (8, 4, 'neigh_op_top_3')
// (8, 5, 'local_g1_3')
// (8, 5, 'lutff_0/in_2')
// (8, 5, 'lutff_3/out')
// (8, 6, 'neigh_op_bot_3')
// (9, 4, 'neigh_op_tnl_3')
// (9, 5, 'neigh_op_lft_3')
// (9, 6, 'neigh_op_bnl_3')

wire n421;
// (7, 4, 'neigh_op_tnr_4')
// (7, 5, 'neigh_op_rgt_4')
// (7, 6, 'neigh_op_bnr_4')
// (8, 4, 'neigh_op_top_4')
// (8, 5, 'lutff_4/out')
// (8, 5, 'sp4_h_r_8')
// (8, 6, 'neigh_op_bot_4')
// (9, 4, 'neigh_op_tnl_4')
// (9, 5, 'neigh_op_lft_4')
// (9, 5, 'sp4_h_r_21')
// (9, 6, 'neigh_op_bnl_4')
// (10, 5, 'sp4_h_r_32')
// (11, 5, 'sp4_h_r_45')
// (11, 6, 'sp4_r_v_b_36')
// (11, 7, 'sp4_r_v_b_25')
// (11, 8, 'sp4_r_v_b_12')
// (11, 9, 'sp4_r_v_b_1')
// (11, 10, 'sp4_r_v_b_36')
// (11, 11, 'local_g0_1')
// (11, 11, 'lutff_3/in_2')
// (11, 11, 'sp4_r_v_b_25')
// (11, 12, 'sp4_r_v_b_12')
// (11, 13, 'sp4_r_v_b_1')
// (12, 5, 'sp4_h_l_45')
// (12, 5, 'sp4_v_t_36')
// (12, 6, 'sp4_v_b_36')
// (12, 7, 'sp4_v_b_25')
// (12, 8, 'sp4_v_b_12')
// (12, 9, 'sp4_v_b_1')
// (12, 9, 'sp4_v_t_36')
// (12, 10, 'sp4_v_b_36')
// (12, 11, 'sp4_v_b_25')
// (12, 12, 'sp4_v_b_12')
// (12, 13, 'sp4_v_b_1')

wire n422;
// (7, 4, 'neigh_op_tnr_5')
// (7, 5, 'neigh_op_rgt_5')
// (7, 6, 'neigh_op_bnr_5')
// (8, 4, 'neigh_op_top_5')
// (8, 5, 'local_g2_5')
// (8, 5, 'lutff_1/in_2')
// (8, 5, 'lutff_5/out')
// (8, 6, 'neigh_op_bot_5')
// (9, 4, 'neigh_op_tnl_5')
// (9, 5, 'neigh_op_lft_5')
// (9, 6, 'neigh_op_bnl_5')

wire n423;
// (7, 4, 'neigh_op_tnr_6')
// (7, 5, 'neigh_op_rgt_6')
// (7, 6, 'neigh_op_bnr_6')
// (8, 4, 'neigh_op_top_6')
// (8, 5, 'local_g2_6')
// (8, 5, 'lutff_0/in_0')
// (8, 5, 'lutff_6/out')
// (8, 6, 'neigh_op_bot_6')
// (9, 4, 'neigh_op_tnl_6')
// (9, 5, 'neigh_op_lft_6')
// (9, 6, 'neigh_op_bnl_6')

wire n424;
// (7, 4, 'neigh_op_tnr_7')
// (7, 5, 'neigh_op_rgt_7')
// (7, 6, 'neigh_op_bnr_7')
// (8, 4, 'neigh_op_top_7')
// (8, 5, 'local_g1_7')
// (8, 5, 'lutff_1/in_1')
// (8, 5, 'lutff_6/in_2')
// (8, 5, 'lutff_7/out')
// (8, 6, 'neigh_op_bot_7')
// (9, 4, 'neigh_op_tnl_7')
// (9, 5, 'neigh_op_lft_7')
// (9, 6, 'neigh_op_bnl_7')

wire n425;
// (7, 5, 'neigh_op_tnr_0')
// (7, 5, 'sp4_r_v_b_45')
// (7, 6, 'neigh_op_rgt_0')
// (7, 6, 'sp4_r_v_b_32')
// (7, 7, 'neigh_op_bnr_0')
// (7, 7, 'sp4_r_v_b_21')
// (7, 8, 'sp4_r_v_b_8')
// (8, 4, 'sp4_v_t_45')
// (8, 5, 'neigh_op_top_0')
// (8, 5, 'sp4_v_b_45')
// (8, 6, 'lutff_0/out')
// (8, 6, 'sp4_v_b_32')
// (8, 7, 'local_g0_0')
// (8, 7, 'local_g1_0')
// (8, 7, 'lutff_2/in_1')
// (8, 7, 'lutff_7/in_1')
// (8, 7, 'neigh_op_bot_0')
// (8, 7, 'sp4_v_b_21')
// (8, 8, 'local_g1_0')
// (8, 8, 'lutff_1/in_2')
// (8, 8, 'sp4_v_b_8')
// (9, 5, 'neigh_op_tnl_0')
// (9, 6, 'neigh_op_lft_0')
// (9, 7, 'neigh_op_bnl_0')

wire n426;
// (7, 5, 'neigh_op_tnr_2')
// (7, 6, 'neigh_op_rgt_2')
// (7, 7, 'neigh_op_bnr_2')
// (8, 5, 'neigh_op_top_2')
// (8, 6, 'lutff_2/out')
// (8, 7, 'local_g0_2')
// (8, 7, 'local_g1_2')
// (8, 7, 'lutff_0/in_3')
// (8, 7, 'lutff_3/in_2')
// (8, 7, 'lutff_4/in_2')
// (8, 7, 'lutff_6/in_2')
// (8, 7, 'neigh_op_bot_2')
// (9, 5, 'neigh_op_tnl_2')
// (9, 6, 'neigh_op_lft_2')
// (9, 7, 'neigh_op_bnl_2')

wire n427;
// (7, 5, 'neigh_op_tnr_3')
// (7, 6, 'neigh_op_rgt_3')
// (7, 7, 'neigh_op_bnr_3')
// (8, 0, 'span12_vert_17')
// (8, 1, 'sp12_v_b_17')
// (8, 2, 'sp12_v_b_14')
// (8, 3, 'sp12_v_b_13')
// (8, 4, 'sp12_v_b_10')
// (8, 5, 'neigh_op_top_3')
// (8, 5, 'sp12_v_b_9')
// (8, 6, 'lutff_3/out')
// (8, 6, 'sp12_v_b_6')
// (8, 7, 'neigh_op_bot_3')
// (8, 7, 'sp12_v_b_5')
// (8, 8, 'local_g2_2')
// (8, 8, 'lutff_3/in_3')
// (8, 8, 'lutff_5/in_1')
// (8, 8, 'sp12_v_b_2')
// (8, 9, 'sp12_v_b_1')
// (9, 5, 'neigh_op_tnl_3')
// (9, 6, 'neigh_op_lft_3')
// (9, 7, 'neigh_op_bnl_3')

wire n428;
// (7, 5, 'neigh_op_tnr_4')
// (7, 6, 'neigh_op_rgt_4')
// (7, 7, 'neigh_op_bnr_4')
// (8, 5, 'neigh_op_top_4')
// (8, 6, 'local_g0_4')
// (8, 6, 'local_g1_4')
// (8, 6, 'lutff_0/in_0')
// (8, 6, 'lutff_1/in_0')
// (8, 6, 'lutff_3/in_0')
// (8, 6, 'lutff_4/out')
// (8, 6, 'lutff_7/in_0')
// (8, 7, 'neigh_op_bot_4')
// (9, 5, 'neigh_op_tnl_4')
// (9, 6, 'neigh_op_lft_4')
// (9, 7, 'neigh_op_bnl_4')

wire n429;
// (7, 5, 'neigh_op_tnr_5')
// (7, 6, 'neigh_op_rgt_5')
// (7, 7, 'neigh_op_bnr_5')
// (8, 5, 'neigh_op_top_5')
// (8, 6, 'lutff_5/out')
// (8, 7, 'local_g0_5')
// (8, 7, 'local_g1_5')
// (8, 7, 'lutff_4/in_0')
// (8, 7, 'lutff_5/in_0')
// (8, 7, 'neigh_op_bot_5')
// (9, 5, 'neigh_op_tnl_5')
// (9, 6, 'neigh_op_lft_5')
// (9, 7, 'neigh_op_bnl_5')

wire n430;
// (7, 5, 'neigh_op_tnr_6')
// (7, 6, 'neigh_op_rgt_6')
// (7, 7, 'neigh_op_bnr_6')
// (8, 5, 'neigh_op_top_6')
// (8, 6, 'local_g1_6')
// (8, 6, 'local_g2_6')
// (8, 6, 'lutff_0/in_1')
// (8, 6, 'lutff_1/in_1')
// (8, 6, 'lutff_3/in_1')
// (8, 6, 'lutff_6/out')
// (8, 6, 'lutff_7/in_1')
// (8, 7, 'neigh_op_bot_6')
// (9, 5, 'neigh_op_tnl_6')
// (9, 6, 'neigh_op_lft_6')
// (9, 7, 'neigh_op_bnl_6')

wire n431;
// (7, 5, 'neigh_op_tnr_7')
// (7, 5, 'sp4_r_v_b_43')
// (7, 6, 'neigh_op_rgt_7')
// (7, 6, 'sp4_r_v_b_30')
// (7, 7, 'neigh_op_bnr_7')
// (7, 7, 'sp4_r_v_b_19')
// (7, 8, 'sp4_r_v_b_6')
// (8, 4, 'sp4_v_t_43')
// (8, 5, 'neigh_op_top_7')
// (8, 5, 'sp4_v_b_43')
// (8, 6, 'lutff_7/out')
// (8, 6, 'sp4_v_b_30')
// (8, 7, 'local_g0_7')
// (8, 7, 'lutff_5/in_2')
// (8, 7, 'neigh_op_bot_7')
// (8, 7, 'sp4_v_b_19')
// (8, 8, 'local_g1_6')
// (8, 8, 'lutff_5/in_2')
// (8, 8, 'sp4_v_b_6')
// (9, 5, 'neigh_op_tnl_7')
// (9, 6, 'neigh_op_lft_7')
// (9, 7, 'neigh_op_bnl_7')

reg n432 = 0;
// (7, 6, 'local_g1_1')
// (7, 6, 'lutff_5/in_3')
// (7, 6, 'sp4_h_r_1')
// (8, 6, 'sp4_h_r_12')
// (9, 6, 'sp4_h_r_25')
// (10, 6, 'neigh_op_tnr_5')
// (10, 6, 'sp4_h_r_36')
// (10, 7, 'neigh_op_rgt_5')
// (10, 7, 'sp4_r_v_b_42')
// (10, 8, 'neigh_op_bnr_5')
// (10, 8, 'sp4_r_v_b_31')
// (10, 9, 'sp4_r_v_b_18')
// (10, 10, 'sp4_r_v_b_7')
// (11, 6, 'local_g0_5')
// (11, 6, 'lutff_0/in_1')
// (11, 6, 'neigh_op_top_5')
// (11, 6, 'sp4_h_l_36')
// (11, 6, 'sp4_v_t_42')
// (11, 7, 'lutff_5/out')
// (11, 7, 'sp4_v_b_42')
// (11, 8, 'neigh_op_bot_5')
// (11, 8, 'sp4_v_b_31')
// (11, 9, 'sp4_v_b_18')
// (11, 10, 'sp4_v_b_7')
// (12, 6, 'neigh_op_tnl_5')
// (12, 7, 'neigh_op_lft_5')
// (12, 8, 'neigh_op_bnl_5')

wire n433;
// (7, 6, 'neigh_op_tnr_0')
// (7, 7, 'neigh_op_rgt_0')
// (7, 8, 'neigh_op_bnr_0')
// (8, 6, 'neigh_op_top_0')
// (8, 7, 'local_g2_0')
// (8, 7, 'lutff_0/out')
// (8, 7, 'lutff_5/in_3')
// (8, 8, 'neigh_op_bot_0')
// (9, 6, 'neigh_op_tnl_0')
// (9, 7, 'neigh_op_lft_0')
// (9, 8, 'neigh_op_bnl_0')

wire n434;
// (7, 6, 'neigh_op_tnr_1')
// (7, 7, 'neigh_op_rgt_1')
// (7, 8, 'neigh_op_bnr_1')
// (8, 6, 'neigh_op_top_1')
// (8, 7, 'local_g0_1')
// (8, 7, 'local_g1_1')
// (8, 7, 'lutff_1/out')
// (8, 7, 'lutff_3/in_0')
// (8, 7, 'lutff_6/in_0')
// (8, 8, 'neigh_op_bot_1')
// (9, 6, 'neigh_op_tnl_1')
// (9, 7, 'neigh_op_lft_1')
// (9, 8, 'neigh_op_bnl_1')

wire n435;
// (7, 6, 'neigh_op_tnr_3')
// (7, 7, 'neigh_op_rgt_3')
// (7, 8, 'neigh_op_bnr_3')
// (8, 6, 'neigh_op_top_3')
// (8, 7, 'local_g0_3')
// (8, 7, 'lutff_2/in_3')
// (8, 7, 'lutff_3/out')
// (8, 7, 'lutff_7/in_2')
// (8, 8, 'neigh_op_bot_3')
// (9, 6, 'neigh_op_tnl_3')
// (9, 7, 'neigh_op_lft_3')
// (9, 8, 'neigh_op_bnl_3')

wire n436;
// (7, 6, 'neigh_op_tnr_4')
// (7, 7, 'neigh_op_rgt_4')
// (7, 8, 'neigh_op_bnr_4')
// (8, 6, 'neigh_op_top_4')
// (8, 7, 'lutff_4/out')
// (8, 8, 'local_g0_4')
// (8, 8, 'local_g1_4')
// (8, 8, 'lutff_4/in_2')
// (8, 8, 'lutff_5/in_0')
// (8, 8, 'lutff_7/in_2')
// (8, 8, 'neigh_op_bot_4')
// (9, 6, 'neigh_op_tnl_4')
// (9, 7, 'neigh_op_lft_4')
// (9, 8, 'neigh_op_bnl_4')

wire n437;
// (7, 6, 'neigh_op_tnr_5')
// (7, 7, 'neigh_op_rgt_5')
// (7, 8, 'neigh_op_bnr_5')
// (8, 0, 'span12_vert_22')
// (8, 1, 'sp12_v_b_22')
// (8, 2, 'sp12_v_b_21')
// (8, 3, 'sp12_v_b_18')
// (8, 4, 'sp12_v_b_17')
// (8, 5, 'sp12_v_b_14')
// (8, 6, 'neigh_op_top_5')
// (8, 6, 'sp12_v_b_13')
// (8, 7, 'lutff_5/out')
// (8, 7, 'sp12_v_b_10')
// (8, 8, 'neigh_op_bot_5')
// (8, 8, 'sp12_v_b_9')
// (8, 9, 'local_g2_6')
// (8, 9, 'lutff_0/in_2')
// (8, 9, 'lutff_1/in_3')
// (8, 9, 'sp12_v_b_6')
// (8, 10, 'sp12_v_b_5')
// (8, 11, 'sp12_v_b_2')
// (8, 12, 'sp12_v_b_1')
// (9, 6, 'neigh_op_tnl_5')
// (9, 7, 'neigh_op_lft_5')
// (9, 8, 'neigh_op_bnl_5')

wire n438;
// (7, 6, 'neigh_op_tnr_6')
// (7, 7, 'neigh_op_rgt_6')
// (7, 8, 'neigh_op_bnr_6')
// (8, 6, 'neigh_op_top_6')
// (8, 7, 'local_g0_6')
// (8, 7, 'lutff_6/out')
// (8, 7, 'lutff_7/in_3')
// (8, 8, 'neigh_op_bot_6')
// (9, 6, 'neigh_op_tnl_6')
// (9, 7, 'neigh_op_lft_6')
// (9, 8, 'neigh_op_bnl_6')

reg n439 = 0;
// (7, 6, 'sp12_h_r_0')
// (8, 5, 'neigh_op_tnr_6')
// (8, 6, 'neigh_op_rgt_6')
// (8, 6, 'sp12_h_r_3')
// (8, 7, 'neigh_op_bnr_6')
// (9, 5, 'neigh_op_top_6')
// (9, 6, 'lutff_6/out')
// (9, 6, 'sp12_h_r_4')
// (9, 7, 'neigh_op_bot_6')
// (10, 5, 'neigh_op_tnl_6')
// (10, 6, 'neigh_op_lft_6')
// (10, 6, 'sp12_h_r_7')
// (10, 7, 'neigh_op_bnl_6')
// (11, 6, 'local_g1_0')
// (11, 6, 'lutff_7/in_0')
// (11, 6, 'sp12_h_r_8')
// (12, 6, 'sp12_h_r_11')
// (13, 6, 'span12_horz_11')

wire n440;
// (7, 6, 'sp4_r_v_b_40')
// (7, 7, 'neigh_op_tnr_0')
// (7, 7, 'sp4_r_v_b_29')
// (7, 8, 'neigh_op_rgt_0')
// (7, 8, 'sp4_r_v_b_16')
// (7, 9, 'neigh_op_bnr_0')
// (7, 9, 'sp4_r_v_b_5')
// (8, 5, 'sp4_r_v_b_36')
// (8, 5, 'sp4_v_t_40')
// (8, 6, 'sp4_r_v_b_25')
// (8, 6, 'sp4_v_b_40')
// (8, 7, 'neigh_op_top_0')
// (8, 7, 'sp4_r_v_b_12')
// (8, 7, 'sp4_v_b_29')
// (8, 8, 'lutff_0/out')
// (8, 8, 'sp4_h_r_0')
// (8, 8, 'sp4_r_v_b_1')
// (8, 8, 'sp4_v_b_16')
// (8, 9, 'local_g0_0')
// (8, 9, 'lutff_6/in_2')
// (8, 9, 'neigh_op_bot_0')
// (8, 9, 'sp4_h_r_5')
// (8, 9, 'sp4_r_v_b_36')
// (8, 9, 'sp4_v_b_5')
// (8, 10, 'sp4_r_v_b_25')
// (8, 11, 'sp4_r_v_b_12')
// (8, 12, 'sp4_r_v_b_1')
// (9, 4, 'sp4_v_t_36')
// (9, 5, 'sp4_v_b_36')
// (9, 6, 'sp4_v_b_25')
// (9, 7, 'neigh_op_tnl_0')
// (9, 7, 'sp4_v_b_12')
// (9, 8, 'neigh_op_lft_0')
// (9, 8, 'sp4_h_r_13')
// (9, 8, 'sp4_v_b_1')
// (9, 8, 'sp4_v_t_36')
// (9, 9, 'neigh_op_bnl_0')
// (9, 9, 'sp4_h_r_16')
// (9, 9, 'sp4_v_b_36')
// (9, 10, 'sp4_v_b_25')
// (9, 11, 'local_g1_4')
// (9, 11, 'lutff_6/in_3')
// (9, 11, 'sp4_v_b_12')
// (9, 12, 'sp4_v_b_1')
// (10, 8, 'sp4_h_r_24')
// (10, 9, 'sp4_h_r_29')
// (11, 8, 'sp4_h_r_37')
// (11, 9, 'local_g2_0')
// (11, 9, 'local_g2_5')
// (11, 9, 'lutff_4/in_3')
// (11, 9, 'lutff_5/in_3')
// (11, 9, 'lutff_6/in_3')
// (11, 9, 'sp4_h_r_40')
// (11, 9, 'sp4_r_v_b_37')
// (11, 10, 'sp4_r_v_b_24')
// (11, 11, 'sp4_r_v_b_13')
// (11, 12, 'sp4_r_v_b_0')
// (12, 8, 'sp4_h_l_37')
// (12, 8, 'sp4_v_t_37')
// (12, 9, 'sp4_h_l_40')
// (12, 9, 'sp4_v_b_37')
// (12, 10, 'sp4_v_b_24')
// (12, 11, 'sp4_v_b_13')
// (12, 12, 'sp4_v_b_0')

wire n441;
// (7, 7, 'neigh_op_tnr_1')
// (7, 8, 'neigh_op_rgt_1')
// (7, 9, 'neigh_op_bnr_1')
// (8, 7, 'neigh_op_top_1')
// (8, 8, 'local_g0_1')
// (8, 8, 'local_g1_1')
// (8, 8, 'lutff_0/in_2')
// (8, 8, 'lutff_1/out')
// (8, 8, 'lutff_2/in_2')
// (8, 8, 'lutff_6/in_1')
// (8, 9, 'neigh_op_bot_1')
// (9, 7, 'neigh_op_tnl_1')
// (9, 8, 'neigh_op_lft_1')
// (9, 9, 'neigh_op_bnl_1')

wire n442;
// (7, 7, 'neigh_op_tnr_2')
// (7, 8, 'neigh_op_rgt_2')
// (7, 8, 'sp4_h_r_9')
// (7, 9, 'neigh_op_bnr_2')
// (8, 7, 'neigh_op_top_2')
// (8, 8, 'lutff_2/out')
// (8, 8, 'sp4_h_r_20')
// (8, 9, 'local_g0_2')
// (8, 9, 'local_g1_2')
// (8, 9, 'lutff_3/in_3')
// (8, 9, 'lutff_4/in_3')
// (8, 9, 'neigh_op_bot_2')
// (9, 7, 'neigh_op_tnl_2')
// (9, 8, 'neigh_op_lft_2')
// (9, 8, 'sp4_h_r_33')
// (9, 9, 'local_g2_2')
// (9, 9, 'lutff_2/in_2')
// (9, 9, 'lutff_5/in_3')
// (9, 9, 'neigh_op_bnl_2')
// (10, 8, 'sp4_h_r_44')
// (10, 9, 'sp4_r_v_b_39')
// (10, 10, 'sp4_r_v_b_26')
// (10, 11, 'sp4_r_v_b_15')
// (10, 12, 'sp4_r_v_b_2')
// (11, 8, 'sp4_h_l_44')
// (11, 8, 'sp4_v_t_39')
// (11, 9, 'local_g2_7')
// (11, 9, 'lutff_2/in_3')
// (11, 9, 'sp4_v_b_39')
// (11, 10, 'sp4_v_b_26')
// (11, 11, 'sp4_v_b_15')
// (11, 12, 'sp4_v_b_2')

wire n443;
// (7, 7, 'neigh_op_tnr_3')
// (7, 8, 'neigh_op_rgt_3')
// (7, 9, 'neigh_op_bnr_3')
// (8, 7, 'neigh_op_top_3')
// (8, 8, 'local_g3_3')
// (8, 8, 'lutff_3/out')
// (8, 8, 'lutff_6/in_2')
// (8, 9, 'neigh_op_bot_3')
// (9, 7, 'neigh_op_tnl_3')
// (9, 8, 'neigh_op_lft_3')
// (9, 9, 'neigh_op_bnl_3')

wire n444;
// (7, 7, 'neigh_op_tnr_4')
// (7, 8, 'neigh_op_rgt_4')
// (7, 9, 'neigh_op_bnr_4')
// (8, 7, 'neigh_op_top_4')
// (8, 8, 'local_g3_4')
// (8, 8, 'lutff_0/in_1')
// (8, 8, 'lutff_4/out')
// (8, 9, 'local_g0_4')
// (8, 9, 'lutff_2/in_2')
// (8, 9, 'neigh_op_bot_4')
// (9, 7, 'neigh_op_tnl_4')
// (9, 8, 'neigh_op_lft_4')
// (9, 9, 'neigh_op_bnl_4')

wire n445;
// (7, 7, 'neigh_op_tnr_5')
// (7, 7, 'sp4_r_v_b_39')
// (7, 8, 'neigh_op_rgt_5')
// (7, 8, 'sp4_r_v_b_26')
// (7, 8, 'sp4_r_v_b_42')
// (7, 9, 'neigh_op_bnr_5')
// (7, 9, 'sp4_r_v_b_15')
// (7, 9, 'sp4_r_v_b_31')
// (7, 10, 'sp4_r_v_b_18')
// (7, 10, 'sp4_r_v_b_2')
// (7, 11, 'sp4_r_v_b_7')
// (8, 6, 'sp4_v_t_39')
// (8, 7, 'neigh_op_top_5')
// (8, 7, 'sp4_h_r_7')
// (8, 7, 'sp4_v_b_39')
// (8, 7, 'sp4_v_t_42')
// (8, 8, 'lutff_5/out')
// (8, 8, 'sp4_v_b_26')
// (8, 8, 'sp4_v_b_42')
// (8, 9, 'local_g0_5')
// (8, 9, 'lutff_0/in_1')
// (8, 9, 'lutff_1/in_2')
// (8, 9, 'neigh_op_bot_5')
// (8, 9, 'sp4_v_b_15')
// (8, 9, 'sp4_v_b_31')
// (8, 10, 'local_g1_2')
// (8, 10, 'lutff_6/in_3')
// (8, 10, 'lutff_7/in_2')
// (8, 10, 'sp4_v_b_18')
// (8, 10, 'sp4_v_b_2')
// (8, 11, 'sp4_v_b_7')
// (9, 7, 'neigh_op_tnl_5')
// (9, 7, 'sp4_h_r_18')
// (9, 8, 'neigh_op_lft_5')
// (9, 9, 'local_g2_5')
// (9, 9, 'local_g3_5')
// (9, 9, 'lutff_2/in_3')
// (9, 9, 'lutff_4/in_3')
// (9, 9, 'lutff_7/in_3')
// (9, 9, 'neigh_op_bnl_5')
// (10, 7, 'sp4_h_r_31')
// (11, 7, 'local_g2_2')
// (11, 7, 'lutff_1/in_3')
// (11, 7, 'sp4_h_r_42')
// (12, 7, 'sp4_h_l_42')

wire n446;
// (7, 7, 'sp4_r_v_b_40')
// (7, 8, 'neigh_op_tnr_0')
// (7, 8, 'sp4_r_v_b_29')
// (7, 9, 'neigh_op_rgt_0')
// (7, 9, 'sp4_r_v_b_16')
// (7, 10, 'neigh_op_bnr_0')
// (7, 10, 'sp4_r_v_b_5')
// (7, 11, 'sp4_r_v_b_36')
// (7, 12, 'sp4_r_v_b_25')
// (7, 13, 'sp4_r_v_b_12')
// (7, 14, 'sp4_r_v_b_1')
// (8, 6, 'sp4_v_t_40')
// (8, 7, 'sp4_v_b_40')
// (8, 8, 'neigh_op_top_0')
// (8, 8, 'sp4_v_b_29')
// (8, 9, 'lutff_0/out')
// (8, 9, 'sp4_v_b_16')
// (8, 10, 'local_g1_5')
// (8, 10, 'lutff_5/in_3')
// (8, 10, 'neigh_op_bot_0')
// (8, 10, 'sp4_v_b_5')
// (8, 10, 'sp4_v_t_36')
// (8, 11, 'sp4_v_b_36')
// (8, 12, 'sp4_v_b_25')
// (8, 13, 'local_g0_4')
// (8, 13, 'local_g1_4')
// (8, 13, 'lutff_1/in_3')
// (8, 13, 'lutff_4/in_3')
// (8, 13, 'lutff_6/in_3')
// (8, 13, 'sp4_v_b_12')
// (8, 14, 'sp4_v_b_1')
// (9, 8, 'neigh_op_tnl_0')
// (9, 9, 'neigh_op_lft_0')
// (9, 10, 'neigh_op_bnl_0')

reg n447 = 0;
// (7, 8, 'neigh_op_tnr_2')
// (7, 9, 'neigh_op_rgt_2')
// (7, 10, 'neigh_op_bnr_2')
// (8, 8, 'neigh_op_top_2')
// (8, 9, 'local_g3_2')
// (8, 9, 'lutff_2/out')
// (8, 9, 'lutff_4/in_1')
// (8, 9, 'lutff_7/in_2')
// (8, 10, 'neigh_op_bot_2')
// (9, 8, 'neigh_op_tnl_2')
// (9, 9, 'neigh_op_lft_2')
// (9, 10, 'neigh_op_bnl_2')

reg n448 = 0;
// (7, 8, 'neigh_op_tnr_3')
// (7, 9, 'local_g3_3')
// (7, 9, 'lutff_0/in_2')
// (7, 9, 'neigh_op_rgt_3')
// (7, 10, 'neigh_op_bnr_3')
// (8, 8, 'neigh_op_top_3')
// (8, 9, 'local_g1_3')
// (8, 9, 'lutff_3/out')
// (8, 9, 'lutff_6/in_0')
// (8, 10, 'neigh_op_bot_3')
// (9, 8, 'neigh_op_tnl_3')
// (9, 9, 'neigh_op_lft_3')
// (9, 10, 'neigh_op_bnl_3')

reg n449 = 0;
// (7, 8, 'neigh_op_tnr_4')
// (7, 9, 'neigh_op_rgt_4')
// (7, 10, 'neigh_op_bnr_4')
// (8, 8, 'neigh_op_top_4')
// (8, 9, 'local_g2_4')
// (8, 9, 'local_g3_4')
// (8, 9, 'lutff_3/in_1')
// (8, 9, 'lutff_4/out')
// (8, 9, 'lutff_5/in_2')
// (8, 10, 'neigh_op_bot_4')
// (9, 8, 'neigh_op_tnl_4')
// (9, 9, 'neigh_op_lft_4')
// (9, 10, 'neigh_op_bnl_4')

reg n450 = 0;
// (7, 8, 'neigh_op_tnr_5')
// (7, 9, 'local_g2_5')
// (7, 9, 'lutff_0/in_1')
// (7, 9, 'neigh_op_rgt_5')
// (7, 10, 'neigh_op_bnr_5')
// (8, 8, 'neigh_op_top_5')
// (8, 9, 'lutff_5/out')
// (8, 10, 'neigh_op_bot_5')
// (9, 8, 'neigh_op_tnl_5')
// (9, 9, 'neigh_op_lft_5')
// (9, 10, 'neigh_op_bnl_5')

reg n451 = 0;
// (7, 8, 'neigh_op_tnr_6')
// (7, 9, 'neigh_op_rgt_6')
// (7, 10, 'neigh_op_bnr_6')
// (8, 8, 'neigh_op_top_6')
// (8, 9, 'local_g1_6')
// (8, 9, 'lutff_2/in_1')
// (8, 9, 'lutff_6/out')
// (8, 10, 'neigh_op_bot_6')
// (9, 8, 'neigh_op_tnl_6')
// (9, 9, 'neigh_op_lft_6')
// (9, 10, 'local_g3_6')
// (9, 10, 'lutff_1/in_0')
// (9, 10, 'neigh_op_bnl_6')

reg n452 = 0;
// (7, 8, 'neigh_op_tnr_7')
// (7, 9, 'neigh_op_rgt_7')
// (7, 10, 'neigh_op_bnr_7')
// (8, 8, 'neigh_op_top_7')
// (8, 9, 'local_g1_7')
// (8, 9, 'lutff_5/in_1')
// (8, 9, 'lutff_7/out')
// (8, 10, 'neigh_op_bot_7')
// (9, 8, 'neigh_op_tnl_7')
// (9, 9, 'neigh_op_lft_7')
// (9, 10, 'neigh_op_bnl_7')

reg n453 = 0;
// (7, 9, 'neigh_op_tnr_0')
// (7, 10, 'local_g3_0')
// (7, 10, 'lutff_1/in_2')
// (7, 10, 'neigh_op_rgt_0')
// (7, 11, 'neigh_op_bnr_0')
// (8, 9, 'neigh_op_top_0')
// (8, 10, 'local_g1_0')
// (8, 10, 'lutff_0/out')
// (8, 10, 'lutff_6/in_1')
// (8, 11, 'neigh_op_bot_0')
// (9, 9, 'neigh_op_tnl_0')
// (9, 10, 'neigh_op_lft_0')
// (9, 11, 'neigh_op_bnl_0')

reg n454 = 0;
// (7, 9, 'neigh_op_tnr_1')
// (7, 10, 'neigh_op_rgt_1')
// (7, 11, 'neigh_op_bnr_1')
// (8, 9, 'neigh_op_top_1')
// (8, 10, 'lutff_1/out')
// (8, 11, 'local_g0_1')
// (8, 11, 'local_g1_1')
// (8, 11, 'lutff_2/in_1')
// (8, 11, 'lutff_6/in_2')
// (8, 11, 'neigh_op_bot_1')
// (9, 9, 'neigh_op_tnl_1')
// (9, 10, 'neigh_op_lft_1')
// (9, 11, 'neigh_op_bnl_1')

reg n455 = 0;
// (7, 9, 'neigh_op_tnr_2')
// (7, 10, 'neigh_op_rgt_2')
// (7, 11, 'neigh_op_bnr_2')
// (8, 9, 'neigh_op_top_2')
// (8, 10, 'local_g3_2')
// (8, 10, 'lutff_0/in_1')
// (8, 10, 'lutff_2/out')
// (8, 10, 'lutff_3/in_2')
// (8, 11, 'neigh_op_bot_2')
// (9, 9, 'neigh_op_tnl_2')
// (9, 10, 'neigh_op_lft_2')
// (9, 11, 'neigh_op_bnl_2')

reg n456 = 0;
// (7, 9, 'neigh_op_tnr_3')
// (7, 10, 'local_g3_3')
// (7, 10, 'lutff_1/in_1')
// (7, 10, 'neigh_op_rgt_3')
// (7, 11, 'neigh_op_bnr_3')
// (8, 9, 'neigh_op_top_3')
// (8, 10, 'lutff_3/out')
// (8, 11, 'neigh_op_bot_3')
// (9, 9, 'neigh_op_tnl_3')
// (9, 10, 'neigh_op_lft_3')
// (9, 11, 'neigh_op_bnl_3')

reg n457 = 0;
// (7, 9, 'neigh_op_tnr_4')
// (7, 10, 'neigh_op_rgt_4')
// (7, 11, 'neigh_op_bnr_4')
// (8, 9, 'neigh_op_top_4')
// (8, 10, 'local_g0_4')
// (8, 10, 'lutff_3/in_1')
// (8, 10, 'lutff_4/out')
// (8, 11, 'neigh_op_bot_4')
// (9, 9, 'neigh_op_tnl_4')
// (9, 10, 'neigh_op_lft_4')
// (9, 11, 'neigh_op_bnl_4')

reg n458 = 0;
// (7, 9, 'neigh_op_tnr_5')
// (7, 10, 'neigh_op_rgt_5')
// (7, 10, 'sp12_h_r_1')
// (7, 11, 'neigh_op_bnr_5')
// (8, 9, 'neigh_op_top_5')
// (8, 10, 'lutff_5/out')
// (8, 10, 'sp12_h_r_2')
// (8, 11, 'neigh_op_bot_5')
// (9, 9, 'neigh_op_tnl_5')
// (9, 10, 'neigh_op_lft_5')
// (9, 10, 'sp12_h_r_5')
// (9, 11, 'neigh_op_bnl_5')
// (10, 10, 'sp12_h_r_6')
// (11, 10, 'local_g0_1')
// (11, 10, 'lutff_1/in_2')
// (11, 10, 'sp12_h_r_9')
// (12, 10, 'sp12_h_r_10')
// (13, 10, 'span12_horz_10')

reg n459 = 0;
// (7, 9, 'neigh_op_tnr_6')
// (7, 10, 'neigh_op_rgt_6')
// (7, 11, 'neigh_op_bnr_6')
// (8, 9, 'neigh_op_top_6')
// (8, 10, 'local_g0_6')
// (8, 10, 'lutff_6/out')
// (8, 10, 'lutff_7/in_1')
// (8, 11, 'neigh_op_bot_6')
// (9, 9, 'neigh_op_tnl_6')
// (9, 10, 'local_g0_6')
// (9, 10, 'lutff_0/in_0')
// (9, 10, 'neigh_op_lft_6')
// (9, 11, 'neigh_op_bnl_6')

reg n460 = 0;
// (7, 9, 'neigh_op_tnr_7')
// (7, 10, 'neigh_op_rgt_7')
// (7, 11, 'neigh_op_bnr_7')
// (8, 9, 'neigh_op_top_7')
// (8, 10, 'local_g0_7')
// (8, 10, 'local_g1_7')
// (8, 10, 'lutff_2/in_1')
// (8, 10, 'lutff_4/in_2')
// (8, 10, 'lutff_7/out')
// (8, 11, 'neigh_op_bot_7')
// (9, 9, 'neigh_op_tnl_7')
// (9, 10, 'neigh_op_lft_7')
// (9, 11, 'neigh_op_bnl_7')

wire \d_out[4] ;
// (7, 9, 'sp12_h_r_0')
// (8, 9, 'sp12_h_r_3')
// (9, 9, 'sp12_h_r_4')
// (10, 8, 'neigh_op_tnr_0')
// (10, 9, 'neigh_op_rgt_0')
// (10, 9, 'sp12_h_r_7')
// (10, 10, 'neigh_op_bnr_0')
// (11, 8, 'neigh_op_top_0')
// (11, 9, 'lutff_0/out')
// (11, 9, 'sp12_h_r_8')
// (11, 10, 'neigh_op_bot_0')
// (12, 8, 'neigh_op_tnl_0')
// (12, 9, 'neigh_op_lft_0')
// (12, 9, 'sp12_h_r_11')
// (12, 10, 'neigh_op_bnl_0')
// (13, 9, 'io_1/D_OUT_0')
// (13, 9, 'io_1/PAD')
// (13, 9, 'local_g0_3')
// (13, 9, 'span12_horz_11')

wire n462;
// (7, 9, 'sp4_r_v_b_40')
// (7, 10, 'local_g0_5')
// (7, 10, 'local_g1_5')
// (7, 10, 'lutff_4/in_1')
// (7, 10, 'lutff_5/in_1')
// (7, 10, 'sp4_r_v_b_29')
// (7, 11, 'sp4_r_v_b_16')
// (7, 12, 'sp4_r_v_b_5')
// (8, 8, 'sp4_v_t_40')
// (8, 9, 'sp4_v_b_40')
// (8, 10, 'sp4_v_b_29')
// (8, 11, 'neigh_op_tnr_0')
// (8, 11, 'sp4_v_b_16')
// (8, 12, 'neigh_op_rgt_0')
// (8, 12, 'sp4_h_r_5')
// (8, 12, 'sp4_v_b_5')
// (8, 13, 'neigh_op_bnr_0')
// (9, 11, 'neigh_op_top_0')
// (9, 12, 'lutff_0/out')
// (9, 12, 'sp4_h_r_16')
// (9, 13, 'neigh_op_bot_0')
// (10, 11, 'neigh_op_tnl_0')
// (10, 12, 'neigh_op_lft_0')
// (10, 12, 'sp4_h_r_29')
// (10, 13, 'neigh_op_bnl_0')
// (11, 12, 'sp4_h_r_40')
// (12, 12, 'sp4_h_l_40')

wire n463;
// (7, 10, 'neigh_op_tnr_0')
// (7, 11, 'local_g3_0')
// (7, 11, 'lutff_2/in_3')
// (7, 11, 'neigh_op_rgt_0')
// (7, 12, 'neigh_op_bnr_0')
// (8, 10, 'neigh_op_top_0')
// (8, 11, 'lutff_0/out')
// (8, 12, 'neigh_op_bot_0')
// (9, 10, 'neigh_op_tnl_0')
// (9, 11, 'neigh_op_lft_0')
// (9, 12, 'neigh_op_bnl_0')

reg n464 = 0;
// (7, 10, 'neigh_op_tnr_1')
// (7, 11, 'local_g3_1')
// (7, 11, 'lutff_2/in_0')
// (7, 11, 'neigh_op_rgt_1')
// (7, 12, 'local_g0_1')
// (7, 12, 'lutff_5/in_0')
// (7, 12, 'neigh_op_bnr_1')
// (8, 10, 'neigh_op_top_1')
// (8, 11, 'local_g2_1')
// (8, 11, 'lutff_1/out')
// (8, 11, 'lutff_7/in_0')
// (8, 12, 'local_g1_1')
// (8, 12, 'lutff_2/in_0')
// (8, 12, 'neigh_op_bot_1')
// (9, 10, 'neigh_op_tnl_1')
// (9, 11, 'neigh_op_lft_1')
// (9, 12, 'neigh_op_bnl_1')

reg n465 = 0;
// (7, 10, 'neigh_op_tnr_2')
// (7, 11, 'local_g3_2')
// (7, 11, 'lutff_4/in_1')
// (7, 11, 'neigh_op_rgt_2')
// (7, 12, 'neigh_op_bnr_2')
// (8, 10, 'neigh_op_top_2')
// (8, 11, 'local_g0_2')
// (8, 11, 'lutff_2/out')
// (8, 11, 'lutff_4/in_2')
// (8, 12, 'neigh_op_bot_2')
// (9, 10, 'neigh_op_tnl_2')
// (9, 11, 'neigh_op_lft_2')
// (9, 12, 'neigh_op_bnl_2')

reg n466 = 0;
// (7, 10, 'neigh_op_tnr_3')
// (7, 11, 'neigh_op_rgt_3')
// (7, 12, 'neigh_op_bnr_3')
// (8, 10, 'neigh_op_top_3')
// (8, 11, 'local_g2_3')
// (8, 11, 'lutff_3/out')
// (8, 11, 'lutff_5/in_0')
// (8, 12, 'neigh_op_bot_3')
// (9, 10, 'neigh_op_tnl_3')
// (9, 11, 'neigh_op_lft_3')
// (9, 12, 'neigh_op_bnl_3')

reg n467 = 0;
// (7, 10, 'neigh_op_tnr_5')
// (7, 11, 'neigh_op_rgt_5')
// (7, 12, 'neigh_op_bnr_5')
// (8, 10, 'neigh_op_top_5')
// (8, 11, 'local_g0_5')
// (8, 11, 'lutff_1/in_0')
// (8, 11, 'lutff_5/out')
// (8, 12, 'neigh_op_bot_5')
// (9, 10, 'neigh_op_tnl_5')
// (9, 11, 'neigh_op_lft_5')
// (9, 12, 'neigh_op_bnl_5')

reg n468 = 0;
// (7, 10, 'neigh_op_tnr_6')
// (7, 11, 'neigh_op_rgt_6')
// (7, 12, 'neigh_op_bnr_6')
// (8, 10, 'neigh_op_top_6')
// (8, 11, 'local_g1_6')
// (8, 11, 'lutff_4/in_1')
// (8, 11, 'lutff_6/out')
// (8, 12, 'neigh_op_bot_6')
// (9, 10, 'neigh_op_tnl_6')
// (9, 11, 'neigh_op_lft_6')
// (9, 12, 'neigh_op_bnl_6')

reg n469 = 0;
// (7, 10, 'neigh_op_tnr_7')
// (7, 11, 'neigh_op_rgt_7')
// (7, 12, 'neigh_op_bnr_7')
// (8, 10, 'neigh_op_top_7')
// (8, 11, 'local_g0_7')
// (8, 11, 'lutff_3/in_0')
// (8, 11, 'lutff_7/out')
// (8, 12, 'neigh_op_bot_7')
// (9, 10, 'neigh_op_tnl_7')
// (9, 11, 'neigh_op_lft_7')
// (9, 12, 'neigh_op_bnl_7')

wire n470;
// (7, 10, 'sp4_r_v_b_37')
// (7, 11, 'local_g0_0')
// (7, 11, 'lutff_1/in_1')
// (7, 11, 'sp4_r_v_b_24')
// (7, 12, 'local_g2_0')
// (7, 12, 'lutff_5/in_1')
// (7, 12, 'neigh_op_tnr_0')
// (7, 12, 'sp4_r_v_b_13')
// (7, 13, 'neigh_op_rgt_0')
// (7, 13, 'sp4_r_v_b_0')
// (7, 14, 'neigh_op_bnr_0')
// (8, 9, 'sp4_v_t_37')
// (8, 10, 'sp4_v_b_37')
// (8, 11, 'sp4_v_b_24')
// (8, 12, 'neigh_op_top_0')
// (8, 12, 'sp4_v_b_13')
// (8, 13, 'lutff_0/out')
// (8, 13, 'sp4_v_b_0')
// (8, 14, 'neigh_op_bot_0')
// (9, 12, 'neigh_op_tnl_0')
// (9, 13, 'neigh_op_lft_0')
// (9, 14, 'neigh_op_bnl_0')

wire n471;
// (7, 11, 'neigh_op_tnr_0')
// (7, 12, 'neigh_op_rgt_0')
// (7, 13, 'neigh_op_bnr_0')
// (8, 10, 'sp4_r_v_b_41')
// (8, 11, 'neigh_op_top_0')
// (8, 11, 'sp4_r_v_b_28')
// (8, 12, 'lutff_0/out')
// (8, 12, 'sp4_h_r_0')
// (8, 12, 'sp4_r_v_b_17')
// (8, 13, 'neigh_op_bot_0')
// (8, 13, 'sp4_r_v_b_4')
// (9, 9, 'sp4_v_t_41')
// (9, 10, 'sp4_v_b_41')
// (9, 11, 'neigh_op_tnl_0')
// (9, 11, 'sp4_v_b_28')
// (9, 12, 'local_g1_1')
// (9, 12, 'lutff_1/in_3')
// (9, 12, 'neigh_op_lft_0')
// (9, 12, 'sp4_h_r_13')
// (9, 12, 'sp4_v_b_17')
// (9, 13, 'neigh_op_bnl_0')
// (9, 13, 'sp4_v_b_4')
// (10, 12, 'sp4_h_r_24')
// (11, 12, 'local_g2_5')
// (11, 12, 'local_g3_5')
// (11, 12, 'lutff_0/in_3')
// (11, 12, 'lutff_7/in_3')
// (11, 12, 'sp4_h_r_37')
// (12, 12, 'sp4_h_l_37')

reg n472 = 0;
// (7, 11, 'neigh_op_tnr_2')
// (7, 12, 'neigh_op_rgt_2')
// (7, 13, 'neigh_op_bnr_2')
// (8, 11, 'neigh_op_top_2')
// (8, 12, 'local_g1_2')
// (8, 12, 'lutff_2/out')
// (8, 12, 'lutff_3/in_0')
// (8, 13, 'neigh_op_bot_2')
// (9, 11, 'neigh_op_tnl_2')
// (9, 12, 'neigh_op_lft_2')
// (9, 13, 'neigh_op_bnl_2')

reg n473 = 0;
// (7, 11, 'neigh_op_tnr_3')
// (7, 12, 'neigh_op_rgt_3')
// (7, 13, 'neigh_op_bnr_3')
// (8, 11, 'neigh_op_top_3')
// (8, 12, 'local_g1_3')
// (8, 12, 'lutff_3/out')
// (8, 12, 'lutff_4/in_0')
// (8, 13, 'neigh_op_bot_3')
// (9, 11, 'neigh_op_tnl_3')
// (9, 12, 'neigh_op_lft_3')
// (9, 13, 'neigh_op_bnl_3')

reg n474 = 0;
// (7, 11, 'neigh_op_tnr_4')
// (7, 12, 'neigh_op_rgt_4')
// (7, 13, 'neigh_op_bnr_4')
// (8, 11, 'neigh_op_top_4')
// (8, 12, 'local_g1_4')
// (8, 12, 'lutff_4/out')
// (8, 12, 'lutff_7/in_0')
// (8, 13, 'neigh_op_bot_4')
// (9, 11, 'neigh_op_tnl_4')
// (9, 12, 'neigh_op_lft_4')
// (9, 13, 'neigh_op_bnl_4')

reg n475 = 0;
// (7, 11, 'neigh_op_tnr_5')
// (7, 11, 'sp4_r_v_b_39')
// (7, 12, 'neigh_op_rgt_5')
// (7, 12, 'sp4_r_v_b_26')
// (7, 13, 'neigh_op_bnr_5')
// (7, 13, 'sp4_r_v_b_15')
// (7, 14, 'sp4_r_v_b_2')
// (8, 10, 'sp4_v_t_39')
// (8, 11, 'local_g2_7')
// (8, 11, 'lutff_0/in_1')
// (8, 11, 'neigh_op_top_5')
// (8, 11, 'sp4_v_b_39')
// (8, 12, 'local_g2_5')
// (8, 12, 'lutff_2/in_1')
// (8, 12, 'lutff_5/out')
// (8, 12, 'sp4_v_b_26')
// (8, 13, 'neigh_op_bot_5')
// (8, 13, 'sp4_v_b_15')
// (8, 14, 'sp4_v_b_2')
// (9, 11, 'neigh_op_tnl_5')
// (9, 12, 'neigh_op_lft_5')
// (9, 13, 'neigh_op_bnl_5')

reg n476 = 0;
// (7, 11, 'neigh_op_tnr_6')
// (7, 12, 'neigh_op_rgt_6')
// (7, 13, 'neigh_op_bnr_6')
// (8, 11, 'neigh_op_top_6')
// (8, 12, 'local_g1_6')
// (8, 12, 'lutff_5/in_0')
// (8, 12, 'lutff_6/out')
// (8, 13, 'neigh_op_bot_6')
// (9, 11, 'neigh_op_tnl_6')
// (9, 12, 'neigh_op_lft_6')
// (9, 13, 'neigh_op_bnl_6')

reg n477 = 0;
// (7, 11, 'neigh_op_tnr_7')
// (7, 12, 'neigh_op_rgt_7')
// (7, 13, 'neigh_op_bnr_7')
// (8, 11, 'local_g1_7')
// (8, 11, 'lutff_0/in_0')
// (8, 11, 'lutff_7/in_1')
// (8, 11, 'neigh_op_top_7')
// (8, 12, 'lutff_7/out')
// (8, 13, 'neigh_op_bot_7')
// (9, 11, 'neigh_op_tnl_7')
// (9, 12, 'neigh_op_lft_7')
// (9, 13, 'neigh_op_bnl_7')

reg n478 = 0;
// (7, 11, 'sp12_h_r_0')
// (8, 10, 'neigh_op_tnr_6')
// (8, 11, 'neigh_op_rgt_6')
// (8, 11, 'sp12_h_r_3')
// (8, 12, 'neigh_op_bnr_6')
// (9, 10, 'neigh_op_top_6')
// (9, 11, 'lutff_6/out')
// (9, 11, 'sp12_h_r_4')
// (9, 12, 'neigh_op_bot_6')
// (10, 10, 'neigh_op_tnl_6')
// (10, 11, 'neigh_op_lft_6')
// (10, 11, 'sp12_h_r_7')
// (10, 12, 'neigh_op_bnl_6')
// (11, 11, 'local_g0_0')
// (11, 11, 'lutff_2/in_2')
// (11, 11, 'sp12_h_r_8')
// (12, 11, 'sp12_h_r_11')
// (13, 11, 'span12_horz_11')

reg n479 = 0;
// (7, 12, 'neigh_op_tnr_1')
// (7, 13, 'neigh_op_rgt_1')
// (7, 14, 'neigh_op_bnr_1')
// (8, 12, 'neigh_op_top_1')
// (8, 13, 'local_g0_1')
// (8, 13, 'local_g1_1')
// (8, 13, 'lutff_1/out')
// (8, 13, 'lutff_2/in_2')
// (8, 13, 'lutff_6/in_1')
// (8, 14, 'neigh_op_bot_1')
// (9, 12, 'neigh_op_tnl_1')
// (9, 13, 'neigh_op_lft_1')
// (9, 14, 'neigh_op_bnl_1')

reg n480 = 0;
// (7, 12, 'neigh_op_tnr_2')
// (7, 13, 'neigh_op_rgt_2')
// (7, 14, 'neigh_op_bnr_2')
// (8, 12, 'neigh_op_top_2')
// (8, 13, 'local_g1_2')
// (8, 13, 'lutff_0/in_1')
// (8, 13, 'lutff_2/out')
// (8, 14, 'neigh_op_bot_2')
// (9, 12, 'neigh_op_tnl_2')
// (9, 13, 'neigh_op_lft_2')
// (9, 14, 'neigh_op_bnl_2')

reg n481 = 0;
// (7, 12, 'neigh_op_tnr_3')
// (7, 13, 'neigh_op_rgt_3')
// (7, 14, 'neigh_op_bnr_3')
// (8, 12, 'neigh_op_top_3')
// (8, 13, 'local_g0_3')
// (8, 13, 'lutff_3/out')
// (8, 13, 'lutff_4/in_1')
// (8, 14, 'local_g0_3')
// (8, 14, 'lutff_3/in_0')
// (8, 14, 'neigh_op_bot_3')
// (9, 12, 'neigh_op_tnl_3')
// (9, 13, 'neigh_op_lft_3')
// (9, 14, 'neigh_op_bnl_3')

reg n482 = 0;
// (7, 12, 'neigh_op_tnr_4')
// (7, 13, 'neigh_op_rgt_4')
// (7, 14, 'neigh_op_bnr_4')
// (8, 12, 'neigh_op_top_4')
// (8, 13, 'local_g2_4')
// (8, 13, 'local_g3_4')
// (8, 13, 'lutff_1/in_1')
// (8, 13, 'lutff_4/out')
// (8, 13, 'lutff_7/in_2')
// (8, 14, 'neigh_op_bot_4')
// (9, 12, 'neigh_op_tnl_4')
// (9, 13, 'neigh_op_lft_4')
// (9, 14, 'neigh_op_bnl_4')

reg n483 = 0;
// (7, 12, 'neigh_op_tnr_6')
// (7, 13, 'neigh_op_rgt_6')
// (7, 14, 'neigh_op_bnr_6')
// (8, 12, 'neigh_op_top_6')
// (8, 13, 'local_g0_6')
// (8, 13, 'lutff_0/in_2')
// (8, 13, 'lutff_3/in_1')
// (8, 13, 'lutff_6/out')
// (8, 14, 'neigh_op_bot_6')
// (9, 12, 'neigh_op_tnl_6')
// (9, 13, 'neigh_op_lft_6')
// (9, 14, 'neigh_op_bnl_6')

reg n484 = 0;
// (7, 12, 'neigh_op_tnr_7')
// (7, 13, 'neigh_op_rgt_7')
// (7, 14, 'neigh_op_bnr_7')
// (8, 12, 'neigh_op_top_7')
// (8, 13, 'local_g0_7')
// (8, 13, 'lutff_2/in_1')
// (8, 13, 'lutff_7/out')
// (8, 14, 'neigh_op_bot_7')
// (9, 12, 'neigh_op_tnl_7')
// (9, 13, 'neigh_op_lft_7')
// (9, 14, 'neigh_op_bnl_7')

reg n485 = 0;
// (7, 12, 'sp12_h_r_0')
// (8, 12, 'sp12_h_r_3')
// (9, 12, 'local_g1_4')
// (9, 12, 'lutff_5/in_2')
// (9, 12, 'sp12_h_r_4')
// (10, 11, 'neigh_op_tnr_0')
// (10, 12, 'neigh_op_rgt_0')
// (10, 12, 'sp12_h_r_7')
// (10, 13, 'neigh_op_bnr_0')
// (11, 11, 'neigh_op_top_0')
// (11, 12, 'local_g0_0')
// (11, 12, 'lutff_0/out')
// (11, 12, 'lutff_3/in_1')
// (11, 12, 'sp12_h_r_8')
// (11, 13, 'neigh_op_bot_0')
// (12, 11, 'neigh_op_tnl_0')
// (12, 12, 'neigh_op_lft_0')
// (12, 12, 'sp12_h_r_11')
// (12, 13, 'neigh_op_bnl_0')
// (13, 12, 'span12_horz_11')

reg n486 = 0;
// (7, 13, 'neigh_op_tnr_3')
// (7, 14, 'neigh_op_rgt_3')
// (7, 15, 'neigh_op_bnr_3')
// (8, 13, 'local_g1_3')
// (8, 13, 'lutff_7/in_1')
// (8, 13, 'neigh_op_top_3')
// (8, 14, 'lutff_3/out')
// (8, 15, 'neigh_op_bot_3')
// (9, 13, 'neigh_op_tnl_3')
// (9, 14, 'neigh_op_lft_3')
// (9, 15, 'neigh_op_bnl_3')

reg n487 = 0;
// (8, 3, 'sp4_h_r_7')
// (9, 3, 'local_g1_2')
// (9, 3, 'lutff_3/in_0')
// (9, 3, 'sp4_h_r_18')
// (10, 2, 'neigh_op_tnr_5')
// (10, 3, 'neigh_op_rgt_5')
// (10, 3, 'sp4_h_r_31')
// (10, 4, 'neigh_op_bnr_5')
// (11, 2, 'neigh_op_top_5')
// (11, 3, 'lutff_5/out')
// (11, 3, 'sp4_h_r_42')
// (11, 4, 'neigh_op_bot_5')
// (12, 2, 'neigh_op_tnl_5')
// (12, 3, 'neigh_op_lft_5')
// (12, 3, 'sp4_h_l_42')
// (12, 4, 'neigh_op_bnl_5')

reg n488 = 0;
// (8, 4, 'neigh_op_tnr_4')
// (8, 5, 'neigh_op_rgt_4')
// (8, 6, 'neigh_op_bnr_4')
// (9, 4, 'neigh_op_top_4')
// (9, 5, 'lutff_4/out')
// (9, 5, 'sp4_h_r_8')
// (9, 6, 'neigh_op_bot_4')
// (10, 4, 'neigh_op_tnl_4')
// (10, 5, 'neigh_op_lft_4')
// (10, 5, 'sp4_h_r_21')
// (10, 6, 'neigh_op_bnl_4')
// (11, 5, 'local_g2_0')
// (11, 5, 'lutff_4/in_0')
// (11, 5, 'sp4_h_r_32')
// (12, 5, 'sp4_h_r_45')
// (13, 5, 'span4_horz_45')

reg n489 = 0;
// (8, 4, 'neigh_op_tnr_7')
// (8, 5, 'neigh_op_rgt_7')
// (8, 6, 'neigh_op_bnr_7')
// (9, 4, 'neigh_op_top_7')
// (9, 5, 'local_g1_7')
// (9, 5, 'lutff_2/in_0')
// (9, 5, 'lutff_7/out')
// (9, 6, 'neigh_op_bot_7')
// (10, 4, 'neigh_op_tnl_7')
// (10, 5, 'neigh_op_lft_7')
// (10, 6, 'neigh_op_bnl_7')

reg n490 = 0;
// (8, 5, 'neigh_op_tnr_3')
// (8, 6, 'neigh_op_rgt_3')
// (8, 6, 'sp4_h_r_11')
// (8, 7, 'neigh_op_bnr_3')
// (9, 5, 'neigh_op_top_3')
// (9, 6, 'lutff_3/out')
// (9, 6, 'sp4_h_r_22')
// (9, 7, 'neigh_op_bot_3')
// (10, 5, 'neigh_op_tnl_3')
// (10, 6, 'neigh_op_lft_3')
// (10, 6, 'sp4_h_r_35')
// (10, 7, 'neigh_op_bnl_3')
// (11, 6, 'local_g3_6')
// (11, 6, 'lutff_1/in_0')
// (11, 6, 'sp4_h_r_46')
// (12, 6, 'sp4_h_l_46')

reg n491 = 0;
// (8, 6, 'neigh_op_tnr_5')
// (8, 6, 'sp4_r_v_b_39')
// (8, 7, 'neigh_op_rgt_5')
// (8, 7, 'sp4_r_v_b_26')
// (8, 8, 'neigh_op_bnr_5')
// (8, 8, 'sp4_r_v_b_15')
// (8, 9, 'sp4_r_v_b_2')
// (9, 5, 'sp4_v_t_39')
// (9, 6, 'neigh_op_top_5')
// (9, 6, 'sp4_v_b_39')
// (9, 7, 'lutff_5/out')
// (9, 7, 'sp4_v_b_26')
// (9, 8, 'neigh_op_bot_5')
// (9, 8, 'sp4_v_b_15')
// (9, 9, 'local_g0_2')
// (9, 9, 'lutff_3/in_1')
// (9, 9, 'sp4_v_b_2')
// (10, 6, 'neigh_op_tnl_5')
// (10, 7, 'neigh_op_lft_5')
// (10, 8, 'neigh_op_bnl_5')

reg n492 = 0;
// (8, 7, 'neigh_op_tnr_0')
// (8, 8, 'neigh_op_rgt_0')
// (8, 9, 'neigh_op_bnr_0')
// (9, 7, 'neigh_op_top_0')
// (9, 8, 'local_g1_0')
// (9, 8, 'lutff_0/out')
// (9, 8, 'lutff_7/in_0')
// (9, 9, 'neigh_op_bot_0')
// (10, 7, 'neigh_op_tnl_0')
// (10, 8, 'neigh_op_lft_0')
// (10, 9, 'neigh_op_bnl_0')

reg n493 = 0;
// (8, 7, 'neigh_op_tnr_1')
// (8, 8, 'neigh_op_rgt_1')
// (8, 9, 'neigh_op_bnr_1')
// (9, 5, 'sp4_r_v_b_38')
// (9, 6, 'local_g0_3')
// (9, 6, 'lutff_6/in_3')
// (9, 6, 'sp4_r_v_b_27')
// (9, 7, 'neigh_op_top_1')
// (9, 7, 'sp4_r_v_b_14')
// (9, 8, 'local_g0_1')
// (9, 8, 'local_g1_1')
// (9, 8, 'lutff_1/out')
// (9, 8, 'lutff_3/in_2')
// (9, 8, 'lutff_5/in_3')
// (9, 8, 'sp4_r_v_b_3')
// (9, 9, 'neigh_op_bot_1')
// (10, 4, 'sp4_v_t_38')
// (10, 5, 'sp4_v_b_38')
// (10, 6, 'sp4_v_b_27')
// (10, 7, 'neigh_op_tnl_1')
// (10, 7, 'sp4_v_b_14')
// (10, 8, 'neigh_op_lft_1')
// (10, 8, 'sp4_h_r_9')
// (10, 8, 'sp4_v_b_3')
// (10, 9, 'neigh_op_bnl_1')
// (11, 8, 'local_g1_4')
// (11, 8, 'lutff_0/in_1')
// (11, 8, 'sp4_h_r_20')
// (12, 8, 'sp4_h_r_33')
// (13, 8, 'span4_horz_33')

reg n494 = 0;
// (8, 7, 'neigh_op_tnr_2')
// (8, 8, 'neigh_op_rgt_2')
// (8, 9, 'neigh_op_bnr_2')
// (9, 7, 'neigh_op_top_2')
// (9, 8, 'local_g0_2')
// (9, 8, 'lutff_2/out')
// (9, 8, 'lutff_4/in_0')
// (9, 9, 'neigh_op_bot_2')
// (10, 7, 'neigh_op_tnl_2')
// (10, 8, 'neigh_op_lft_2')
// (10, 9, 'neigh_op_bnl_2')

reg n495 = 0;
// (8, 7, 'neigh_op_tnr_3')
// (8, 8, 'neigh_op_rgt_3')
// (8, 9, 'neigh_op_bnr_3')
// (9, 7, 'neigh_op_top_3')
// (9, 8, 'local_g1_3')
// (9, 8, 'lutff_0/in_0')
// (9, 8, 'lutff_3/out')
// (9, 9, 'neigh_op_bot_3')
// (10, 7, 'neigh_op_tnl_3')
// (10, 8, 'neigh_op_lft_3')
// (10, 9, 'neigh_op_bnl_3')

reg n496 = 0;
// (8, 7, 'neigh_op_tnr_4')
// (8, 8, 'neigh_op_rgt_4')
// (8, 9, 'neigh_op_bnr_4')
// (9, 7, 'neigh_op_top_4')
// (9, 8, 'local_g2_4')
// (9, 8, 'lutff_3/in_3')
// (9, 8, 'lutff_4/out')
// (9, 9, 'neigh_op_bot_4')
// (10, 7, 'neigh_op_tnl_4')
// (10, 8, 'neigh_op_lft_4')
// (10, 9, 'neigh_op_bnl_4')

reg n497 = 0;
// (8, 7, 'neigh_op_tnr_7')
// (8, 8, 'neigh_op_rgt_7')
// (8, 9, 'neigh_op_bnr_7')
// (9, 7, 'neigh_op_top_7')
// (9, 8, 'local_g0_7')
// (9, 8, 'lutff_1/in_0')
// (9, 8, 'lutff_7/out')
// (9, 9, 'neigh_op_bot_7')
// (10, 7, 'neigh_op_tnl_7')
// (10, 8, 'neigh_op_lft_7')
// (10, 9, 'neigh_op_bnl_7')

reg n498 = 0;
// (8, 8, 'neigh_op_tnr_2')
// (8, 9, 'neigh_op_rgt_2')
// (8, 10, 'neigh_op_bnr_2')
// (9, 8, 'neigh_op_top_2')
// (9, 9, 'local_g1_2')
// (9, 9, 'lutff_2/out')
// (9, 9, 'lutff_3/in_2')
// (9, 9, 'lutff_4/in_1')
// (9, 10, 'neigh_op_bot_2')
// (10, 8, 'neigh_op_tnl_2')
// (10, 9, 'neigh_op_lft_2')
// (10, 10, 'neigh_op_bnl_2')

reg n499 = 0;
// (8, 8, 'neigh_op_tnr_3')
// (8, 9, 'neigh_op_rgt_3')
// (8, 10, 'neigh_op_bnr_3')
// (9, 8, 'neigh_op_top_3')
// (9, 9, 'local_g0_3')
// (9, 9, 'lutff_3/out')
// (9, 9, 'lutff_6/in_1')
// (9, 10, 'neigh_op_bot_3')
// (10, 8, 'neigh_op_tnl_3')
// (10, 9, 'neigh_op_lft_3')
// (10, 10, 'neigh_op_bnl_3')

reg n500 = 0;
// (8, 8, 'neigh_op_tnr_4')
// (8, 9, 'neigh_op_rgt_4')
// (8, 10, 'neigh_op_bnr_4')
// (9, 8, 'neigh_op_top_4')
// (9, 9, 'local_g0_4')
// (9, 9, 'lutff_4/out')
// (9, 9, 'lutff_6/in_2')
// (9, 9, 'lutff_7/in_1')
// (9, 10, 'neigh_op_bot_4')
// (10, 8, 'neigh_op_tnl_4')
// (10, 9, 'neigh_op_lft_4')
// (10, 10, 'neigh_op_bnl_4')

reg n501 = 0;
// (8, 8, 'neigh_op_tnr_5')
// (8, 9, 'neigh_op_rgt_5')
// (8, 10, 'neigh_op_bnr_5')
// (9, 6, 'sp4_r_v_b_46')
// (9, 7, 'local_g2_3')
// (9, 7, 'lutff_5/in_0')
// (9, 7, 'sp4_r_v_b_35')
// (9, 8, 'neigh_op_top_5')
// (9, 8, 'sp4_r_v_b_22')
// (9, 9, 'local_g0_5')
// (9, 9, 'lutff_2/in_1')
// (9, 9, 'lutff_5/out')
// (9, 9, 'sp4_r_v_b_11')
// (9, 10, 'neigh_op_bot_5')
// (10, 5, 'sp4_v_t_46')
// (10, 6, 'sp4_v_b_46')
// (10, 7, 'sp4_v_b_35')
// (10, 8, 'neigh_op_tnl_5')
// (10, 8, 'sp4_v_b_22')
// (10, 9, 'neigh_op_lft_5')
// (10, 9, 'sp4_v_b_11')
// (10, 10, 'neigh_op_bnl_5')

reg n502 = 0;
// (8, 8, 'neigh_op_tnr_6')
// (8, 9, 'neigh_op_rgt_6')
// (8, 10, 'neigh_op_bnr_6')
// (9, 8, 'neigh_op_top_6')
// (9, 9, 'local_g0_6')
// (9, 9, 'lutff_1/in_1')
// (9, 9, 'lutff_6/out')
// (9, 10, 'neigh_op_bot_6')
// (10, 8, 'neigh_op_tnl_6')
// (10, 9, 'neigh_op_lft_6')
// (10, 10, 'neigh_op_bnl_6')

reg n503 = 0;
// (8, 8, 'neigh_op_tnr_7')
// (8, 9, 'neigh_op_rgt_7')
// (8, 10, 'neigh_op_bnr_7')
// (9, 8, 'neigh_op_top_7')
// (9, 9, 'local_g0_7')
// (9, 9, 'local_g1_7')
// (9, 9, 'lutff_1/in_2')
// (9, 9, 'lutff_5/in_1')
// (9, 9, 'lutff_7/out')
// (9, 10, 'neigh_op_bot_7')
// (10, 8, 'neigh_op_tnl_7')
// (10, 9, 'neigh_op_lft_7')
// (10, 10, 'neigh_op_bnl_7')

reg n504 = 0;
// (8, 9, 'local_g3_1')
// (8, 9, 'lutff_7/in_1')
// (8, 9, 'neigh_op_tnr_1')
// (8, 10, 'neigh_op_rgt_1')
// (8, 11, 'neigh_op_bnr_1')
// (9, 9, 'neigh_op_top_1')
// (9, 10, 'lutff_1/out')
// (9, 11, 'neigh_op_bot_1')
// (10, 9, 'neigh_op_tnl_1')
// (10, 10, 'neigh_op_lft_1')
// (10, 11, 'neigh_op_bnl_1')

reg n505 = 0;
// (8, 9, 'neigh_op_tnr_0')
// (8, 10, 'local_g3_0')
// (8, 10, 'lutff_4/in_1')
// (8, 10, 'neigh_op_rgt_0')
// (8, 11, 'neigh_op_bnr_0')
// (9, 9, 'neigh_op_top_0')
// (9, 10, 'lutff_0/out')
// (9, 11, 'neigh_op_bot_0')
// (10, 9, 'neigh_op_tnl_0')
// (10, 10, 'neigh_op_lft_0')
// (10, 11, 'neigh_op_bnl_0')

reg n506 = 0;
// (8, 9, 'sp4_h_r_11')
// (9, 9, 'local_g1_6')
// (9, 9, 'lutff_0/in_1')
// (9, 9, 'sp4_h_r_22')
// (10, 8, 'neigh_op_tnr_7')
// (10, 9, 'neigh_op_rgt_7')
// (10, 9, 'sp4_h_r_35')
// (10, 10, 'neigh_op_bnr_7')
// (11, 8, 'neigh_op_top_7')
// (11, 9, 'lutff_7/out')
// (11, 9, 'sp4_h_r_46')
// (11, 10, 'neigh_op_bot_7')
// (12, 8, 'neigh_op_tnl_7')
// (12, 9, 'neigh_op_lft_7')
// (12, 9, 'sp4_h_l_46')
// (12, 10, 'neigh_op_bnl_7')

reg n507 = 0;
// (8, 10, 'neigh_op_tnr_1')
// (8, 11, 'neigh_op_rgt_1')
// (8, 12, 'neigh_op_bnr_1')
// (9, 10, 'neigh_op_top_1')
// (9, 11, 'local_g1_1')
// (9, 11, 'lutff_1/out')
// (9, 11, 'lutff_2/in_0')
// (9, 12, 'neigh_op_bot_1')
// (10, 10, 'neigh_op_tnl_1')
// (10, 11, 'neigh_op_lft_1')
// (10, 12, 'neigh_op_bnl_1')

reg n508 = 0;
// (8, 10, 'neigh_op_tnr_2')
// (8, 11, 'neigh_op_rgt_2')
// (8, 12, 'neigh_op_bnr_2')
// (9, 10, 'neigh_op_top_2')
// (9, 11, 'local_g1_2')
// (9, 11, 'lutff_2/out')
// (9, 11, 'lutff_3/in_0')
// (9, 12, 'neigh_op_bot_2')
// (10, 10, 'neigh_op_tnl_2')
// (10, 11, 'neigh_op_lft_2')
// (10, 12, 'neigh_op_bnl_2')

reg n509 = 0;
// (8, 10, 'neigh_op_tnr_5')
// (8, 11, 'neigh_op_rgt_5')
// (8, 12, 'neigh_op_bnr_5')
// (9, 4, 'sp12_v_t_22')
// (9, 5, 'sp12_v_b_22')
// (9, 6, 'sp12_v_b_21')
// (9, 7, 'sp12_v_b_18')
// (9, 8, 'local_g3_1')
// (9, 8, 'lutff_2/in_0')
// (9, 8, 'sp12_v_b_17')
// (9, 9, 'sp12_v_b_14')
// (9, 10, 'neigh_op_top_5')
// (9, 10, 'sp12_v_b_13')
// (9, 11, 'lutff_5/out')
// (9, 11, 'sp12_v_b_10')
// (9, 12, 'neigh_op_bot_5')
// (9, 12, 'sp12_v_b_9')
// (9, 13, 'sp12_v_b_6')
// (9, 14, 'sp12_v_b_5')
// (9, 15, 'sp12_v_b_2')
// (9, 16, 'sp12_v_b_1')
// (10, 10, 'neigh_op_tnl_5')
// (10, 11, 'neigh_op_lft_5')
// (10, 12, 'neigh_op_bnl_5')

reg n510 = 0;
// (8, 10, 'neigh_op_tnr_7')
// (8, 11, 'neigh_op_rgt_7')
// (8, 12, 'neigh_op_bnr_7')
// (9, 10, 'neigh_op_top_7')
// (9, 11, 'local_g0_7')
// (9, 11, 'lutff_1/in_0')
// (9, 11, 'lutff_7/out')
// (9, 12, 'neigh_op_bot_7')
// (10, 10, 'neigh_op_tnl_7')
// (10, 11, 'neigh_op_lft_7')
// (10, 12, 'neigh_op_bnl_7')

reg n511 = 0;
// (8, 11, 'neigh_op_tnr_1')
// (8, 12, 'neigh_op_rgt_1')
// (8, 12, 'sp4_h_r_7')
// (8, 13, 'neigh_op_bnr_1')
// (9, 11, 'neigh_op_top_1')
// (9, 12, 'lutff_1/out')
// (9, 12, 'sp4_h_r_18')
// (9, 13, 'neigh_op_bot_1')
// (10, 11, 'neigh_op_tnl_1')
// (10, 12, 'neigh_op_lft_1')
// (10, 12, 'sp4_h_r_31')
// (10, 13, 'neigh_op_bnl_1')
// (11, 9, 'sp4_r_v_b_42')
// (11, 10, 'sp4_r_v_b_31')
// (11, 11, 'local_g3_2')
// (11, 11, 'lutff_5/in_0')
// (11, 11, 'sp4_r_v_b_18')
// (11, 12, 'local_g2_2')
// (11, 12, 'lutff_7/in_1')
// (11, 12, 'sp4_h_r_42')
// (11, 12, 'sp4_r_v_b_7')
// (12, 8, 'sp4_v_t_42')
// (12, 9, 'sp4_v_b_42')
// (12, 10, 'sp4_v_b_31')
// (12, 11, 'sp4_v_b_18')
// (12, 12, 'sp4_h_l_42')
// (12, 12, 'sp4_v_b_7')

reg n512 = 0;
// (8, 11, 'neigh_op_tnr_2')
// (8, 12, 'local_g2_2')
// (8, 12, 'lutff_1/in_1')
// (8, 12, 'neigh_op_rgt_2')
// (8, 13, 'neigh_op_bnr_2')
// (9, 11, 'neigh_op_top_2')
// (9, 12, 'lutff_2/out')
// (9, 13, 'neigh_op_bot_2')
// (10, 11, 'neigh_op_tnl_2')
// (10, 12, 'neigh_op_lft_2')
// (10, 13, 'neigh_op_bnl_2')

reg n513 = 0;
// (8, 11, 'neigh_op_tnr_3')
// (8, 12, 'neigh_op_rgt_3')
// (8, 13, 'neigh_op_bnr_3')
// (9, 11, 'neigh_op_top_3')
// (9, 12, 'local_g2_3')
// (9, 12, 'lutff_3/out')
// (9, 12, 'lutff_4/in_1')
// (9, 13, 'neigh_op_bot_3')
// (10, 11, 'neigh_op_tnl_3')
// (10, 12, 'neigh_op_lft_3')
// (10, 13, 'neigh_op_bnl_3')

reg n514 = 0;
// (8, 11, 'neigh_op_tnr_4')
// (8, 12, 'neigh_op_rgt_4')
// (8, 13, 'neigh_op_bnr_4')
// (9, 11, 'neigh_op_top_4')
// (9, 12, 'local_g3_4')
// (9, 12, 'lutff_0/in_1')
// (9, 12, 'lutff_4/out')
// (9, 13, 'neigh_op_bot_4')
// (10, 11, 'neigh_op_tnl_4')
// (10, 12, 'neigh_op_lft_4')
// (10, 13, 'neigh_op_bnl_4')

reg n515 = 0;
// (8, 11, 'neigh_op_tnr_5')
// (8, 12, 'neigh_op_rgt_5')
// (8, 13, 'neigh_op_bnr_5')
// (9, 11, 'neigh_op_top_5')
// (9, 12, 'local_g0_5')
// (9, 12, 'lutff_2/in_1')
// (9, 12, 'lutff_5/out')
// (9, 13, 'neigh_op_bot_5')
// (10, 11, 'neigh_op_tnl_5')
// (10, 12, 'neigh_op_lft_5')
// (10, 13, 'neigh_op_bnl_5')

reg n516 = 0;
// (8, 11, 'neigh_op_tnr_6')
// (8, 12, 'neigh_op_rgt_6')
// (8, 12, 'sp4_h_r_1')
// (8, 13, 'neigh_op_bnr_6')
// (9, 11, 'neigh_op_top_6')
// (9, 12, 'lutff_6/out')
// (9, 12, 'sp4_h_r_12')
// (9, 13, 'neigh_op_bot_6')
// (10, 11, 'neigh_op_tnl_6')
// (10, 12, 'neigh_op_lft_6')
// (10, 12, 'sp4_h_r_25')
// (10, 13, 'neigh_op_bnl_6')
// (11, 9, 'sp4_r_v_b_36')
// (11, 10, 'sp4_r_v_b_25')
// (11, 11, 'sp4_r_v_b_12')
// (11, 12, 'local_g2_4')
// (11, 12, 'lutff_0/in_2')
// (11, 12, 'sp4_h_r_36')
// (11, 12, 'sp4_r_v_b_1')
// (12, 8, 'sp4_v_t_36')
// (12, 9, 'sp4_v_b_36')
// (12, 10, 'sp4_v_b_25')
// (12, 11, 'sp4_v_b_12')
// (12, 12, 'local_g0_1')
// (12, 12, 'lutff_7/in_0')
// (12, 12, 'sp4_h_l_36')
// (12, 12, 'sp4_v_b_1')

reg n517 = 0;
// (8, 11, 'neigh_op_tnr_7')
// (8, 12, 'neigh_op_rgt_7')
// (8, 13, 'neigh_op_bnr_7')
// (9, 11, 'neigh_op_top_7')
// (9, 12, 'local_g1_7')
// (9, 12, 'lutff_0/in_2')
// (9, 12, 'lutff_1/in_1')
// (9, 12, 'lutff_7/out')
// (9, 13, 'neigh_op_bot_7')
// (10, 11, 'neigh_op_tnl_7')
// (10, 12, 'neigh_op_lft_7')
// (10, 13, 'neigh_op_bnl_7')

wire n518;
// (8, 11, 'sp4_h_r_3')
// (9, 11, 'local_g0_6')
// (9, 11, 'local_g1_6')
// (9, 11, 'lutff_6/in_2')
// (9, 11, 'lutff_7/in_2')
// (9, 11, 'sp4_h_r_14')
// (10, 10, 'neigh_op_tnr_3')
// (10, 11, 'neigh_op_rgt_3')
// (10, 11, 'sp4_h_r_27')
// (10, 12, 'neigh_op_bnr_3')
// (11, 10, 'local_g1_3')
// (11, 10, 'lutff_6/in_0')
// (11, 10, 'neigh_op_top_3')
// (11, 11, 'lutff_3/out')
// (11, 11, 'sp4_h_r_38')
// (11, 12, 'neigh_op_bot_3')
// (12, 10, 'neigh_op_tnl_3')
// (12, 11, 'neigh_op_lft_3')
// (12, 11, 'sp4_h_l_38')
// (12, 12, 'neigh_op_bnl_3')

reg n519 = 0;
// (8, 12, 'neigh_op_tnr_2')
// (8, 13, 'neigh_op_rgt_2')
// (8, 14, 'neigh_op_bnr_2')
// (9, 12, 'neigh_op_top_2')
// (9, 13, 'local_g1_2')
// (9, 13, 'lutff_2/out')
// (9, 13, 'lutff_5/in_0')
// (9, 14, 'neigh_op_bot_2')
// (10, 12, 'neigh_op_tnl_2')
// (10, 13, 'neigh_op_lft_2')
// (10, 14, 'neigh_op_bnl_2')

reg n520 = 0;
// (8, 12, 'neigh_op_tnr_3')
// (8, 13, 'neigh_op_rgt_3')
// (8, 14, 'neigh_op_bnr_3')
// (9, 12, 'neigh_op_top_3')
// (9, 13, 'lutff_3/out')
// (9, 14, 'local_g1_3')
// (9, 14, 'lutff_4/in_0')
// (9, 14, 'neigh_op_bot_3')
// (10, 12, 'neigh_op_tnl_3')
// (10, 13, 'neigh_op_lft_3')
// (10, 14, 'neigh_op_bnl_3')

reg n521 = 0;
// (8, 12, 'neigh_op_tnr_6')
// (8, 13, 'neigh_op_rgt_6')
// (8, 14, 'neigh_op_bnr_6')
// (9, 12, 'neigh_op_top_6')
// (9, 13, 'local_g1_6')
// (9, 13, 'lutff_3/in_0')
// (9, 13, 'lutff_6/out')
// (9, 14, 'neigh_op_bot_6')
// (10, 12, 'neigh_op_tnl_6')
// (10, 13, 'neigh_op_lft_6')
// (10, 14, 'neigh_op_bnl_6')

reg n522 = 0;
// (8, 12, 'neigh_op_tnr_7')
// (8, 13, 'neigh_op_rgt_7')
// (8, 14, 'neigh_op_bnr_7')
// (9, 12, 'neigh_op_top_7')
// (9, 13, 'local_g1_7')
// (9, 13, 'lutff_6/in_0')
// (9, 13, 'lutff_7/out')
// (9, 14, 'neigh_op_bot_7')
// (10, 12, 'neigh_op_tnl_7')
// (10, 13, 'neigh_op_lft_7')
// (10, 14, 'neigh_op_bnl_7')

reg n523 = 0;
// (8, 12, 'sp4_h_r_3')
// (9, 12, 'local_g0_6')
// (9, 12, 'lutff_2/in_2')
// (9, 12, 'sp4_h_r_14')
// (10, 11, 'neigh_op_tnr_3')
// (10, 12, 'neigh_op_rgt_3')
// (10, 12, 'sp4_h_r_27')
// (10, 13, 'neigh_op_bnr_3')
// (11, 11, 'neigh_op_top_3')
// (11, 12, 'local_g1_3')
// (11, 12, 'lutff_1/in_1')
// (11, 12, 'lutff_3/out')
// (11, 12, 'sp4_h_r_38')
// (11, 13, 'neigh_op_bot_3')
// (12, 11, 'neigh_op_tnl_3')
// (12, 12, 'neigh_op_lft_3')
// (12, 12, 'sp4_h_l_38')
// (12, 13, 'neigh_op_bnl_3')

reg n524 = 0;
// (8, 12, 'sp4_r_v_b_45')
// (8, 13, 'sp4_r_v_b_32')
// (8, 14, 'sp4_r_v_b_21')
// (8, 15, 'sp4_r_v_b_8')
// (9, 11, 'sp4_h_r_2')
// (9, 11, 'sp4_v_t_45')
// (9, 12, 'local_g3_5')
// (9, 12, 'lutff_3/in_1')
// (9, 12, 'sp4_v_b_45')
// (9, 13, 'sp4_v_b_32')
// (9, 14, 'sp4_v_b_21')
// (9, 15, 'sp4_v_b_8')
// (10, 10, 'neigh_op_tnr_5')
// (10, 11, 'neigh_op_rgt_5')
// (10, 11, 'sp4_h_r_15')
// (10, 12, 'neigh_op_bnr_5')
// (11, 10, 'neigh_op_top_5')
// (11, 11, 'lutff_5/out')
// (11, 11, 'sp4_h_r_26')
// (11, 12, 'neigh_op_bot_5')
// (12, 10, 'neigh_op_tnl_5')
// (12, 11, 'neigh_op_lft_5')
// (12, 11, 'sp4_h_r_39')
// (12, 12, 'neigh_op_bnl_5')
// (13, 11, 'span4_horz_39')

reg n525 = 0;
// (8, 13, 'neigh_op_tnr_1')
// (8, 14, 'neigh_op_rgt_1')
// (8, 15, 'neigh_op_bnr_1')
// (9, 13, 'neigh_op_top_1')
// (9, 14, 'local_g1_1')
// (9, 14, 'lutff_1/out')
// (9, 14, 'lutff_6/in_0')
// (9, 15, 'neigh_op_bot_1')
// (10, 13, 'neigh_op_tnl_1')
// (10, 14, 'neigh_op_lft_1')
// (10, 15, 'neigh_op_bnl_1')

reg n526 = 0;
// (8, 13, 'neigh_op_tnr_3')
// (8, 14, 'neigh_op_rgt_3')
// (8, 15, 'neigh_op_bnr_3')
// (9, 13, 'neigh_op_top_3')
// (9, 14, 'local_g0_3')
// (9, 14, 'lutff_3/out')
// (9, 14, 'lutff_5/in_0')
// (9, 15, 'neigh_op_bot_3')
// (10, 13, 'neigh_op_tnl_3')
// (10, 14, 'neigh_op_lft_3')
// (10, 15, 'neigh_op_bnl_3')

reg n527 = 0;
// (8, 13, 'neigh_op_tnr_4')
// (8, 14, 'neigh_op_rgt_4')
// (8, 15, 'neigh_op_bnr_4')
// (9, 13, 'neigh_op_top_4')
// (9, 14, 'local_g1_4')
// (9, 14, 'lutff_1/in_0')
// (9, 14, 'lutff_4/out')
// (9, 15, 'neigh_op_bot_4')
// (10, 13, 'neigh_op_tnl_4')
// (10, 14, 'neigh_op_lft_4')
// (10, 15, 'neigh_op_bnl_4')

reg n528 = 0;
// (8, 13, 'neigh_op_tnr_5')
// (8, 14, 'neigh_op_rgt_5')
// (8, 15, 'neigh_op_bnr_5')
// (9, 7, 'sp12_v_t_22')
// (9, 8, 'sp12_v_b_22')
// (9, 9, 'sp12_v_b_21')
// (9, 10, 'sp12_v_b_18')
// (9, 11, 'local_g3_1')
// (9, 11, 'lutff_7/in_3')
// (9, 11, 'sp12_v_b_17')
// (9, 12, 'sp12_v_b_14')
// (9, 13, 'neigh_op_top_5')
// (9, 13, 'sp12_v_b_13')
// (9, 14, 'lutff_5/out')
// (9, 14, 'sp12_v_b_10')
// (9, 15, 'neigh_op_bot_5')
// (9, 15, 'sp12_v_b_9')
// (9, 16, 'sp12_v_b_6')
// (9, 17, 'span12_vert_5')
// (10, 13, 'neigh_op_tnl_5')
// (10, 14, 'neigh_op_lft_5')
// (10, 15, 'neigh_op_bnl_5')

reg n529 = 0;
// (8, 13, 'neigh_op_tnr_6')
// (8, 14, 'neigh_op_rgt_6')
// (8, 15, 'neigh_op_bnr_6')
// (9, 13, 'neigh_op_top_6')
// (9, 14, 'local_g1_6')
// (9, 14, 'lutff_3/in_0')
// (9, 14, 'lutff_6/out')
// (9, 15, 'neigh_op_bot_6')
// (10, 13, 'neigh_op_tnl_6')
// (10, 14, 'neigh_op_lft_6')
// (10, 15, 'neigh_op_bnl_6')

reg n530 = 0;
// (8, 13, 'sp12_h_r_1')
// (9, 13, 'local_g0_2')
// (9, 13, 'lutff_2/in_0')
// (9, 13, 'sp12_h_r_2')
// (10, 12, 'neigh_op_tnr_7')
// (10, 13, 'neigh_op_rgt_7')
// (10, 13, 'sp12_h_r_5')
// (10, 14, 'neigh_op_bnr_7')
// (11, 12, 'neigh_op_top_7')
// (11, 13, 'lutff_7/out')
// (11, 13, 'sp12_h_r_6')
// (11, 14, 'neigh_op_bot_7')
// (12, 12, 'neigh_op_tnl_7')
// (12, 13, 'neigh_op_lft_7')
// (12, 13, 'sp12_h_r_9')
// (12, 14, 'neigh_op_bnl_7')
// (13, 13, 'span12_horz_9')

reg n531 = 0;
// (9, 5, 'local_g1_2')
// (9, 5, 'lutff_7/in_0')
// (9, 5, 'sp4_h_r_10')
// (10, 4, 'neigh_op_tnr_1')
// (10, 5, 'neigh_op_rgt_1')
// (10, 5, 'sp4_h_r_23')
// (10, 6, 'neigh_op_bnr_1')
// (11, 4, 'neigh_op_top_1')
// (11, 5, 'lutff_1/out')
// (11, 5, 'sp4_h_r_34')
// (11, 6, 'neigh_op_bot_1')
// (12, 4, 'neigh_op_tnl_1')
// (12, 5, 'neigh_op_lft_1')
// (12, 5, 'sp4_h_r_47')
// (12, 6, 'neigh_op_bnl_1')
// (13, 5, 'span4_horz_47')

reg n532 = 0;
// (9, 12, 'local_g1_3')
// (9, 12, 'lutff_5/in_1')
// (9, 12, 'sp4_h_r_11')
// (10, 12, 'sp4_h_r_22')
// (11, 11, 'neigh_op_tnr_7')
// (11, 12, 'neigh_op_rgt_7')
// (11, 12, 'sp4_h_r_35')
// (11, 13, 'neigh_op_bnr_7')
// (12, 11, 'neigh_op_top_7')
// (12, 12, 'lutff_7/out')
// (12, 12, 'sp4_h_r_46')
// (12, 13, 'neigh_op_bot_7')
// (13, 11, 'logic_op_tnl_7')
// (13, 12, 'logic_op_lft_7')
// (13, 12, 'span4_horz_46')
// (13, 13, 'logic_op_bnl_7')

reg n533 = 0;
// (10, 3, 'neigh_op_tnr_5')
// (10, 4, 'neigh_op_rgt_5')
// (10, 5, 'neigh_op_bnr_5')
// (11, 3, 'local_g0_5')
// (11, 3, 'lutff_5/in_0')
// (11, 3, 'neigh_op_top_5')
// (11, 4, 'lutff_5/out')
// (11, 5, 'neigh_op_bot_5')
// (12, 3, 'neigh_op_tnl_5')
// (12, 4, 'neigh_op_lft_5')
// (12, 5, 'neigh_op_bnl_5')

reg n534 = 0;
// (10, 4, 'neigh_op_tnr_4')
// (10, 5, 'neigh_op_rgt_4')
// (10, 6, 'neigh_op_bnr_4')
// (11, 4, 'neigh_op_top_4')
// (11, 5, 'local_g0_4')
// (11, 5, 'lutff_1/in_3')
// (11, 5, 'lutff_4/out')
// (11, 6, 'neigh_op_bot_4')
// (12, 4, 'neigh_op_tnl_4')
// (12, 5, 'neigh_op_lft_4')
// (12, 6, 'neigh_op_bnl_4')

reg n535 = 0;
// (10, 5, 'neigh_op_tnr_1')
// (10, 6, 'neigh_op_rgt_1')
// (10, 7, 'neigh_op_bnr_1')
// (11, 5, 'neigh_op_top_1')
// (11, 6, 'local_g0_1')
// (11, 6, 'lutff_1/out')
// (11, 6, 'lutff_5/in_0')
// (11, 7, 'neigh_op_bot_1')
// (12, 5, 'neigh_op_tnl_1')
// (12, 6, 'neigh_op_lft_1')
// (12, 7, 'neigh_op_bnl_1')

reg n536 = 0;
// (10, 5, 'neigh_op_tnr_7')
// (10, 6, 'neigh_op_rgt_7')
// (10, 7, 'neigh_op_bnr_7')
// (11, 5, 'local_g0_7')
// (11, 5, 'lutff_3/in_0')
// (11, 5, 'neigh_op_top_7')
// (11, 6, 'lutff_7/out')
// (11, 7, 'neigh_op_bot_7')
// (12, 5, 'neigh_op_tnl_7')
// (12, 6, 'neigh_op_lft_7')
// (12, 7, 'neigh_op_bnl_7')

reg n537 = 0;
// (10, 6, 'neigh_op_tnr_0')
// (10, 7, 'neigh_op_rgt_0')
// (10, 8, 'neigh_op_bnr_0')
// (11, 6, 'neigh_op_top_0')
// (11, 6, 'sp4_r_v_b_44')
// (11, 7, 'local_g0_2')
// (11, 7, 'lutff_0/out')
// (11, 7, 'lutff_7/in_3')
// (11, 7, 'sp4_r_v_b_33')
// (11, 8, 'neigh_op_bot_0')
// (11, 8, 'sp4_r_v_b_20')
// (11, 9, 'sp4_r_v_b_9')
// (12, 5, 'sp4_v_t_44')
// (12, 6, 'neigh_op_tnl_0')
// (12, 6, 'sp4_v_b_44')
// (12, 7, 'neigh_op_lft_0')
// (12, 7, 'sp4_v_b_33')
// (12, 8, 'neigh_op_bnl_0')
// (12, 8, 'sp4_v_b_20')
// (12, 9, 'sp4_v_b_9')

reg n538 = 0;
// (10, 6, 'neigh_op_tnr_1')
// (10, 7, 'neigh_op_rgt_1')
// (10, 8, 'neigh_op_bnr_1')
// (11, 6, 'local_g1_1')
// (11, 6, 'lutff_0/in_2')
// (11, 6, 'neigh_op_top_1')
// (11, 7, 'lutff_1/out')
// (11, 8, 'neigh_op_bot_1')
// (12, 6, 'neigh_op_tnl_1')
// (12, 7, 'neigh_op_lft_1')
// (12, 8, 'neigh_op_bnl_1')

reg n539 = 0;
// (10, 6, 'neigh_op_tnr_2')
// (10, 7, 'neigh_op_rgt_2')
// (10, 8, 'neigh_op_bnr_2')
// (11, 6, 'neigh_op_top_2')
// (11, 7, 'local_g1_2')
// (11, 7, 'lutff_2/out')
// (11, 7, 'lutff_5/in_0')
// (11, 8, 'neigh_op_bot_2')
// (12, 6, 'neigh_op_tnl_2')
// (12, 7, 'neigh_op_lft_2')
// (12, 8, 'neigh_op_bnl_2')

reg n540 = 0;
// (10, 6, 'neigh_op_tnr_4')
// (10, 7, 'neigh_op_rgt_4')
// (10, 8, 'neigh_op_bnr_4')
// (11, 6, 'neigh_op_top_4')
// (11, 7, 'local_g0_4')
// (11, 7, 'lutff_2/in_0')
// (11, 7, 'lutff_4/out')
// (11, 8, 'neigh_op_bot_4')
// (12, 6, 'neigh_op_tnl_4')
// (12, 7, 'neigh_op_lft_4')
// (12, 8, 'neigh_op_bnl_4')

reg n541 = 0;
// (10, 6, 'neigh_op_tnr_7')
// (10, 7, 'neigh_op_rgt_7')
// (10, 8, 'neigh_op_bnr_7')
// (11, 6, 'neigh_op_top_7')
// (11, 7, 'local_g1_7')
// (11, 7, 'lutff_4/in_0')
// (11, 7, 'lutff_7/out')
// (11, 8, 'neigh_op_bot_7')
// (12, 6, 'neigh_op_tnl_7')
// (12, 7, 'neigh_op_lft_7')
// (12, 8, 'neigh_op_bnl_7')

wire \d_out[1] ;
// (10, 7, 'neigh_op_tnr_0')
// (10, 8, 'neigh_op_rgt_0')
// (10, 9, 'neigh_op_bnr_0')
// (11, 7, 'neigh_op_top_0')
// (11, 8, 'lutff_0/out')
// (11, 8, 'sp4_h_r_0')
// (11, 9, 'neigh_op_bot_0')
// (12, 7, 'neigh_op_tnl_0')
// (12, 8, 'neigh_op_lft_0')
// (12, 8, 'sp4_h_r_13')
// (12, 9, 'neigh_op_bnl_0')
// (13, 8, 'span4_horz_13')
// (13, 8, 'span4_vert_t_14')
// (13, 9, 'span4_vert_b_14')
// (13, 10, 'span4_vert_b_10')
// (13, 11, 'span4_vert_b_6')
// (13, 12, 'io_0/D_OUT_0')
// (13, 12, 'io_0/PAD')
// (13, 12, 'local_g0_2')
// (13, 12, 'span4_vert_b_2')

wire \d_out[0] ;
// (10, 7, 'neigh_op_tnr_1')
// (10, 8, 'neigh_op_rgt_1')
// (10, 8, 'sp4_h_r_7')
// (10, 9, 'neigh_op_bnr_1')
// (11, 7, 'neigh_op_top_1')
// (11, 8, 'lutff_1/out')
// (11, 8, 'sp4_h_r_18')
// (11, 9, 'neigh_op_bot_1')
// (12, 7, 'neigh_op_tnl_1')
// (12, 8, 'neigh_op_lft_1')
// (12, 8, 'sp4_h_r_31')
// (12, 9, 'neigh_op_bnl_1')
// (13, 8, 'span4_horz_31')
// (13, 8, 'span4_vert_t_13')
// (13, 9, 'span4_vert_b_13')
// (13, 10, 'span4_vert_b_9')
// (13, 11, 'span4_vert_b_5')
// (13, 12, 'io_1/D_OUT_0')
// (13, 12, 'io_1/PAD')
// (13, 12, 'local_g0_1')
// (13, 12, 'span4_vert_b_1')

reg n544 = 0;
// (10, 7, 'neigh_op_tnr_2')
// (10, 8, 'neigh_op_rgt_2')
// (10, 9, 'neigh_op_bnr_2')
// (11, 7, 'neigh_op_top_2')
// (11, 8, 'local_g1_2')
// (11, 8, 'lutff_1/in_2')
// (11, 8, 'lutff_2/out')
// (11, 9, 'neigh_op_bot_2')
// (12, 7, 'neigh_op_tnl_2')
// (12, 8, 'neigh_op_lft_2')
// (12, 9, 'neigh_op_bnl_2')

reg n545 = 0;
// (10, 7, 'neigh_op_tnr_7')
// (10, 8, 'neigh_op_rgt_7')
// (10, 9, 'neigh_op_bnr_7')
// (11, 7, 'neigh_op_top_7')
// (11, 8, 'local_g0_7')
// (11, 8, 'lutff_3/in_0')
// (11, 8, 'lutff_7/out')
// (11, 9, 'neigh_op_bot_7')
// (12, 7, 'neigh_op_tnl_7')
// (12, 8, 'neigh_op_lft_7')
// (12, 9, 'neigh_op_bnl_7')

reg n546 = 0;
// (10, 8, 'neigh_op_tnr_1')
// (10, 9, 'neigh_op_rgt_1')
// (10, 10, 'neigh_op_bnr_1')
// (11, 8, 'neigh_op_top_1')
// (11, 9, 'local_g0_1')
// (11, 9, 'lutff_1/out')
// (11, 9, 'lutff_4/in_1')
// (11, 10, 'neigh_op_bot_1')
// (12, 8, 'neigh_op_tnl_1')
// (12, 9, 'local_g0_1')
// (12, 9, 'lutff_5/in_0')
// (12, 9, 'neigh_op_lft_1')
// (12, 10, 'neigh_op_bnl_1')

reg n547 = 0;
// (10, 8, 'neigh_op_tnr_2')
// (10, 9, 'neigh_op_rgt_2')
// (10, 10, 'neigh_op_bnr_2')
// (11, 8, 'neigh_op_top_2')
// (11, 9, 'local_g0_2')
// (11, 9, 'lutff_0/in_2')
// (11, 9, 'lutff_2/out')
// (11, 10, 'neigh_op_bot_2')
// (12, 8, 'neigh_op_tnl_2')
// (12, 9, 'neigh_op_lft_2')
// (12, 10, 'neigh_op_bnl_2')

reg n548 = 0;
// (10, 8, 'neigh_op_tnr_3')
// (10, 9, 'neigh_op_rgt_3')
// (10, 10, 'neigh_op_bnr_3')
// (11, 8, 'neigh_op_top_3')
// (11, 9, 'local_g1_3')
// (11, 9, 'lutff_3/out')
// (11, 9, 'lutff_7/in_1')
// (11, 10, 'neigh_op_bot_3')
// (12, 8, 'neigh_op_tnl_3')
// (12, 9, 'neigh_op_lft_3')
// (12, 10, 'neigh_op_bnl_3')

reg n549 = 0;
// (10, 8, 'neigh_op_tnr_4')
// (10, 9, 'neigh_op_rgt_4')
// (10, 10, 'neigh_op_bnr_4')
// (11, 8, 'neigh_op_top_4')
// (11, 9, 'local_g0_4')
// (11, 9, 'local_g1_4')
// (11, 9, 'lutff_3/in_2')
// (11, 9, 'lutff_4/out')
// (11, 9, 'lutff_5/in_1')
// (11, 10, 'neigh_op_bot_4')
// (12, 8, 'neigh_op_tnl_4')
// (12, 9, 'neigh_op_lft_4')
// (12, 10, 'neigh_op_bnl_4')

reg n550 = 0;
// (10, 8, 'neigh_op_tnr_5')
// (10, 9, 'neigh_op_rgt_5')
// (10, 10, 'neigh_op_bnr_5')
// (11, 8, 'neigh_op_top_5')
// (11, 9, 'local_g0_5')
// (11, 9, 'lutff_5/out')
// (11, 9, 'lutff_6/in_1')
// (11, 9, 'lutff_7/in_2')
// (11, 10, 'neigh_op_bot_5')
// (12, 8, 'neigh_op_tnl_5')
// (12, 9, 'neigh_op_lft_5')
// (12, 10, 'neigh_op_bnl_5')

wire \d_out[2] ;
// (10, 9, 'neigh_op_tnr_1')
// (10, 10, 'neigh_op_rgt_1')
// (10, 10, 'sp4_h_r_7')
// (10, 11, 'neigh_op_bnr_1')
// (11, 9, 'neigh_op_top_1')
// (11, 10, 'lutff_1/out')
// (11, 10, 'sp4_h_r_18')
// (11, 11, 'neigh_op_bot_1')
// (12, 9, 'neigh_op_tnl_1')
// (12, 10, 'neigh_op_lft_1')
// (12, 10, 'sp4_h_r_31')
// (12, 11, 'neigh_op_bnl_1')
// (13, 10, 'span4_horz_31')
// (13, 10, 'span4_vert_t_13')
// (13, 11, 'io_1/D_OUT_0')
// (13, 11, 'io_1/PAD')
// (13, 11, 'local_g0_5')
// (13, 11, 'span4_vert_b_13')
// (13, 12, 'span4_vert_b_9')
// (13, 13, 'span4_vert_b_5')
// (13, 14, 'span4_vert_b_1')

reg n552 = 0;
// (10, 9, 'neigh_op_tnr_6')
// (10, 10, 'neigh_op_rgt_6')
// (10, 11, 'neigh_op_bnr_6')
// (11, 8, 'local_g2_5')
// (11, 8, 'lutff_7/in_0')
// (11, 8, 'sp4_r_v_b_37')
// (11, 9, 'neigh_op_top_6')
// (11, 9, 'sp4_r_v_b_24')
// (11, 10, 'lutff_6/out')
// (11, 10, 'sp4_r_v_b_13')
// (11, 11, 'neigh_op_bot_6')
// (11, 11, 'sp4_r_v_b_0')
// (12, 7, 'sp4_v_t_37')
// (12, 8, 'sp4_v_b_37')
// (12, 9, 'neigh_op_tnl_6')
// (12, 9, 'sp4_v_b_24')
// (12, 10, 'neigh_op_lft_6')
// (12, 10, 'sp4_v_b_13')
// (12, 11, 'neigh_op_bnl_6')
// (12, 11, 'sp4_v_b_0')

wire \d_out[3] ;
// (10, 10, 'neigh_op_tnr_2')
// (10, 11, 'neigh_op_rgt_2')
// (10, 11, 'sp4_h_r_9')
// (10, 12, 'neigh_op_bnr_2')
// (11, 10, 'neigh_op_top_2')
// (11, 11, 'lutff_2/out')
// (11, 11, 'sp4_h_r_20')
// (11, 12, 'neigh_op_bot_2')
// (12, 10, 'neigh_op_tnl_2')
// (12, 11, 'neigh_op_lft_2')
// (12, 11, 'sp4_h_r_33')
// (12, 12, 'neigh_op_bnl_2')
// (13, 11, 'io_0/D_OUT_0')
// (13, 11, 'io_0/PAD')
// (13, 11, 'local_g1_1')
// (13, 11, 'span4_horz_33')

reg n554 = 0;
// (11, 8, 'neigh_op_tnr_5')
// (11, 9, 'local_g3_5')
// (11, 9, 'lutff_3/in_1')
// (11, 9, 'neigh_op_rgt_5')
// (11, 10, 'neigh_op_bnr_5')
// (12, 8, 'neigh_op_top_5')
// (12, 9, 'lutff_5/out')
// (12, 10, 'neigh_op_bot_5')
// (13, 8, 'logic_op_tnl_5')
// (13, 9, 'logic_op_lft_5')
// (13, 10, 'logic_op_bnl_5')

reg n555 = 0;
// (11, 9, 'neigh_op_tnr_0')
// (11, 10, 'neigh_op_rgt_0')
// (11, 11, 'neigh_op_bnr_0')
// (12, 9, 'neigh_op_top_0')
// (12, 10, 'local_g1_0')
// (12, 10, 'lutff_0/out')
// (12, 10, 'lutff_1/in_0')
// (12, 11, 'neigh_op_bot_0')
// (13, 9, 'logic_op_tnl_0')
// (13, 10, 'logic_op_lft_0')
// (13, 11, 'logic_op_bnl_0')

reg n556 = 0;
// (11, 9, 'neigh_op_tnr_1')
// (11, 10, 'neigh_op_rgt_1')
// (11, 11, 'neigh_op_bnr_1')
// (12, 9, 'neigh_op_top_1')
// (12, 10, 'lutff_1/out')
// (12, 11, 'local_g1_1')
// (12, 11, 'lutff_2/in_0')
// (12, 11, 'neigh_op_bot_1')
// (13, 9, 'logic_op_tnl_1')
// (13, 10, 'logic_op_lft_1')
// (13, 11, 'logic_op_bnl_1')

reg n557 = 0;
// (11, 10, 'neigh_op_tnr_2')
// (11, 11, 'neigh_op_rgt_2')
// (11, 12, 'neigh_op_bnr_2')
// (12, 10, 'neigh_op_top_2')
// (12, 11, 'local_g1_2')
// (12, 11, 'lutff_2/out')
// (12, 11, 'lutff_5/in_0')
// (12, 12, 'neigh_op_bot_2')
// (13, 10, 'logic_op_tnl_2')
// (13, 11, 'logic_op_lft_2')
// (13, 12, 'logic_op_bnl_2')

reg n558 = 0;
// (11, 10, 'neigh_op_tnr_5')
// (11, 11, 'neigh_op_rgt_5')
// (11, 12, 'neigh_op_bnr_5')
// (12, 10, 'neigh_op_top_5')
// (12, 11, 'local_g0_5')
// (12, 11, 'lutff_5/out')
// (12, 11, 'lutff_7/in_0')
// (12, 12, 'neigh_op_bot_5')
// (13, 10, 'logic_op_tnl_5')
// (13, 11, 'logic_op_lft_5')
// (13, 12, 'logic_op_bnl_5')

wire n559;
// (2, 5, 'lutff_0/cout')

wire n560;
// (1, 3, 'lutff_0/cout')

wire n561;
// (5, 12, 'lutff_6/lout')

wire n562;
// (9, 12, 'lutff_1/lout')

wire n563;
// (2, 8, 'lutff_3/lout')

wire n564;
// (6, 8, 'lutff_4/lout')

wire n565;
// (4, 8, 'lutff_5/lout')

wire n566;
// (8, 8, 'lutff_6/lout')

wire n567;
// (7, 4, 'lutff_4/lout')

wire n568;
// (1, 7, 'lutff_4/lout')

wire n569;
// (7, 13, 'lutff_0/lout')

wire n570;
// (9, 13, 'lutff_2/lout')

wire n571;
// (5, 5, 'lutff_3/lout')

wire n572;
// (7, 5, 'lutff_5/lout')

wire n573;
// (4, 12, 'lutff_2/lout')

wire n574;
// (8, 12, 'lutff_3/lout')

wire n575;
// (9, 5, 'lutff_7/lout')

wire n576;
// (6, 4, 'lutff_6/lout')

wire n577;
// (5, 9, 'lutff_0/lout')

wire n578;
// (7, 9, 'lutff_2/lout')

wire n579;
// (9, 9, 'lutff_4/lout')

wire n580;
// (5, 8, 'lutff_4/lout')

wire n581;
// (7, 8, 'lutff_6/lout')

wire n582;
// (1, 3, 'lutff_2/lout')

wire n583;
// (8, 11, 'lutff_7/lout')

wire n584;
// (11, 6, 'lutff_5/lout')

wire n585;
// (5, 12, 'lutff_1/lout')

wire n586;
// (7, 12, 'lutff_3/lout')

wire n587;
// (9, 12, 'lutff_5/lout')

wire n588;
// (8, 8, 'lutff_1/lout')

wire n589;
// (7, 13, 'lutff_4/lout')

wire n590;
// (7, 5, 'lutff_0/lout')

wire n591;
// (9, 13, 'lutff_6/lout')

wire n592;
// (5, 5, 'lutff_7/lout')

wire n593;
// (9, 5, 'lutff_2/lout')

wire n594;
// (12, 9, 'lutff_5/lout')

wire n595;
// (4, 12, 'lutff_6/lout')

wire n596;
// (8, 4, 'lutff_3/lout')

wire n597;
// (6, 7, 'lutff_3/lout')

wire n598;
// (8, 7, 'lutff_5/lout')

wire n599;
// (7, 8, 'lutff_1/lout')

wire n600;
// (9, 8, 'lutff_3/lout')

wire n601;
// (5, 11, 'lutff_4/lout')

wire n602;
// (7, 11, 'lutff_6/lout')

wire n603;
// (4, 7, 'lutff_3/lout')

wire n604;
// (6, 11, 'lutff_0/lout')

wire n605;
// (11, 6, 'lutff_0/lout')

wire n606;
// (8, 11, 'lutff_2/lout')

wire n607;
// (11, 9, 'lutff_5/lout')

wire n608;
// (9, 12, 'lutff_0/lout')

wire n609;
// (6, 8, 'lutff_3/lout')

wire n610;
// (7, 12, 'lutff_7/lout')

wire n611;
// (4, 8, 'lutff_4/lout')

wire n612;
// (7, 4, 'lutff_3/lout')

wire n613;
// (8, 8, 'lutff_5/lout')

wire n614;
// (11, 10, 'lutff_6/lout')

wire n615;
// (8, 3, 'lutff_3/lout')

wire n616;
// (6, 6, 'lutff_6/lout')

wire n617;
// (8, 7, 'lutff_0/lout')

wire n618;
// (6, 7, 'lutff_7/lout')

wire n619;
// (11, 13, 'lutff_7/lout')

wire n620;
// (11, 5, 'lutff_3/lout')

wire n621;
// (1, 6, 'lutff_7/lout')

wire n622;
// (5, 8, 'lutff_3/lout')

wire n623;
// (7, 8, 'lutff_5/lout')

wire n624;
// (7, 11, 'lutff_1/lout')

wire n625;
// (9, 8, 'lutff_7/lout')

wire n626;
// (1, 3, 'lutff_1/out')

wire n627;
// (1, 3, 'lutff_1/lout')

wire n628;
// (6, 11, 'lutff_4/lout')

wire n629;
// (11, 6, 'lutff_4/lout')

wire n630;
// (8, 11, 'lutff_6/lout')

wire n631;
// (11, 9, 'lutff_0/lout')

wire n632;
// (5, 12, 'lutff_0/lout')

wire n633;
// (7, 12, 'lutff_2/lout')

wire n634;
// (9, 12, 'lutff_4/lout')

wire n635;
// (5, 4, 'lutff_5/lout')

wire n636;
// (7, 4, 'lutff_7/lout')

wire n637;
// (11, 10, 'lutff_1/lout')

wire n638;
// (6, 6, 'lutff_1/lout')

wire n639;
// (8, 3, 'lutff_7/lout')

wire n640;
// (4, 11, 'lutff_0/lout')

wire n641;
// (2, 3, 'lutff_3/lout')

wire n642;
// (2, 14, 'lutff_3/lout')

wire n643;
// (4, 3, 'lutff_5/lout')

wire n644;
// (6, 7, 'lutff_2/lout')

wire n645;
// (8, 7, 'lutff_4/lout')

wire n646;
// (7, 8, 'lutff_0/lout')

wire n647;
// (5, 8, 'lutff_7/lout')

wire n648;
// (9, 8, 'lutff_2/lout')

wire n649;
// (5, 11, 'lutff_3/lout')

wire n650;
// (7, 11, 'lutff_5/lout')

wire n651;
// (4, 7, 'lutff_2/lout')

wire n652;
// (8, 11, 'lutff_1/lout')

wire n653;
// (6, 10, 'lutff_3/lout')

wire n654;
// (11, 9, 'lutff_4/lout')

wire n655;
// (8, 10, 'lutff_5/lout')

wire n656;
// (5, 4, 'lutff_0/lout')

wire n657;
// (7, 4, 'lutff_2/lout')

wire n658;
// (9, 11, 'lutff_3/lout')

wire n659;
// (2, 10, 'lutff_1/lout')

wire n660;
// (7, 3, 'lutff_6/lout')

wire n661;
// (6, 3, 'lutff_0/lout')

wire n662;
// (8, 3, 'lutff_2/lout')

wire n663;
// (2, 2, 'lutff_6/lout')

wire n664;
// (6, 6, 'lutff_5/lout')

wire n665;
// (9, 4, 'lutff_0/lout')

wire n666;
// (7, 15, 'lutff_7/lout')

wire n667;
// (4, 11, 'lutff_4/lout')

wire n668;
// (7, 7, 'lutff_3/lout')

wire n669;
// (4, 3, 'lutff_0/lout')

wire n670;
// (9, 7, 'lutff_5/lout')

wire n671;
// (2, 3, 'lutff_7/lout')

wire n672;
// (5, 8, 'lutff_2/lout')

wire n673;
// (7, 8, 'lutff_4/lout')

wire n674;
// (7, 11, 'lutff_0/lout')

wire n675;
// (5, 11, 'lutff_7/lout')

wire n676;
// (8, 10, 'lutff_0/lout')

wire n677;
// (6, 10, 'lutff_7/lout')

wire n678;
// (6, 13, 'lutff_3/lout')

wire n679;
// (8, 2, 'lutff_5/lout')

wire n680;
// (9, 11, 'lutff_7/lout')

wire n681;
// (7, 3, 'lutff_1/lout')

wire n682;
// (9, 3, 'lutff_3/lout')

wire n683;
// (5, 6, 'lutff_4/lout')

wire n684;
// (2, 2, 'lutff_1/lout')

wire n685;
// (6, 3, 'lutff_4/lout')

wire n686;
// (4, 10, 'lutff_7/lout')

wire n687;
// (8, 3, 'lutff_6/lout')

wire n688;
// (11, 12, 'lutff_0/lout')

wire n689;
// (7, 15, 'lutff_2/lout')

wire n690;
// (11, 4, 'lutff_5/lout')

wire n691;
// (5, 7, 'lutff_5/lout')

wire n692;
// (2, 3, 'lutff_2/lout')

wire n693;
// (7, 7, 'lutff_7/lout')

wire n694;
// (8, 6, 'lutff_7/lout')

wire n695;
// (6, 9, 'lutff_1/lout')

wire n696;
// (2, 6, 'lutff_3/lout')

wire n697;
// (5, 14, 'lutff_4/lout')

wire n698;
// (6, 10, 'lutff_2/lout')

wire n699;
// (7, 14, 'lutff_6/lout')

wire n700;
// (8, 10, 'lutff_4/lout')

wire n701;
// (8, 2, 'lutff_0/lout')

wire n702;
// (6, 13, 'lutff_7/lout')

wire n703;
// (6, 2, 'lutff_7/lout')

wire n704;
// (11, 8, 'lutff_7/lout')

wire n705;
// (9, 11, 'lutff_2/lout')

wire n706;
// (2, 10, 'lutff_0/lout')

wire n707;
// (7, 3, 'lutff_5/lout')

wire n708;
// (4, 10, 'lutff_2/lout')

wire n709;
// (9, 3, 'lutff_7/lout')

wire n710;
// (8, 3, 'lutff_1/lout')

wire n711;
// (4, 2, 'lutff_7/lout')

wire n712;
// (7, 7, 'lutff_2/lout')

wire n713;
// (5, 10, 'lutff_2/lout')

wire n714;
// (7, 10, 'lutff_4/lout')

wire n715;
// (11, 5, 'lutff_1/lout')

wire n716;
// (8, 6, 'lutff_2/lout')

wire n717;
// (6, 9, 'lutff_5/lout')

wire n718;
// (4, 9, 'lutff_6/lout')

wire n719;
// (8, 9, 'lutff_7/lout')

wire n720;
// (4, 6, 'lutff_0/lout')

wire n721;
// (7, 14, 'lutff_1/lout')

wire n722;
// (2, 6, 'lutff_7/lout')

wire n723;
// (9, 14, 'lutff_3/lout')

wire n724;
// (6, 10, 'lutff_6/lout')

wire n725;
// (6, 2, 'lutff_2/lout')

wire n726;
// (6, 13, 'lutff_2/lout')

wire n727;
// (11, 8, 'lutff_2/lout')

wire n728;
// (8, 2, 'lutff_4/lout')

wire n729;
// (7, 3, 'lutff_0/lout')

wire n730;
// (9, 11, 'lutff_6/lout')

wire n731;
// (2, 10, 'lutff_4/lout')

wire n732;
// (5, 6, 'lutff_3/lout')

wire n733;
// (4, 10, 'lutff_6/lout')

wire n734;
// (8, 13, 'lutff_0/lout')

wire n735;
// (6, 5, 'lutff_3/lout')

wire n736;
// (8, 5, 'lutff_5/lout')

wire n737;
// (5, 10, 'lutff_6/lout')

wire n738;
// (9, 10, 'lutff_1/lout')

wire n739;
// (5, 13, 'lutff_2/lout')

wire n740;
// (6, 9, 'lutff_0/lout')

wire n741;
// (8, 6, 'lutff_6/lout')

wire n742;
// (4, 9, 'lutff_1/lout')

wire n743;
// (8, 9, 'lutff_2/lout')

wire n744;
// (7, 2, 'lutff_4/lout')

wire n745;
// (11, 7, 'lutff_5/lout')

wire n746;
// (2, 6, 'lutff_2/lout')

wire n747;
// (4, 6, 'lutff_4/lout')

wire n748;
// (7, 14, 'lutff_5/lout')

wire n749;
// (6, 10, 'lutff_1/lout')

wire n750;
// (8, 10, 'lutff_3/lout')

wire n751;
// (6, 13, 'lutff_6/lout')

wire n752;
// (9, 11, 'lutff_1/lout')

wire n753;
// (7, 3, 'lutff_4/lout')

wire n754;
// (4, 10, 'lutff_1/lout')

wire n755;
// (5, 6, 'lutff_7/lout')

wire n756;
// (2, 2, 'lutff_4/lout')

wire n757;
// (7, 6, 'lutff_6/lout')

wire n758;
// (11, 12, 'lutff_3/lout')

wire n759;
// (8, 13, 'lutff_4/lout')

wire n760;
// (8, 5, 'lutff_0/lout')

wire n761;
// (2, 5, 'lutff_6/lout')

wire n762;
// (6, 5, 'lutff_7/lout')

wire n763;
// (5, 10, 'lutff_1/lout')

wire n764;
// (7, 10, 'lutff_3/lout')

wire n765;
// (8, 6, 'lutff_1/lout')

wire n766;
// (2, 9, 'lutff_3/lout')

wire n767;
// (6, 9, 'lutff_4/lout')

wire n768;
// (4, 9, 'lutff_5/lout')

wire n769;
// (8, 9, 'lutff_6/lout')

wire n770;
// (11, 7, 'lutff_0/lout')

wire n771;
// (7, 14, 'lutff_0/lout')

wire n772;
// (2, 6, 'lutff_6/lout')

wire n773;
// (11, 8, 'lutff_1/lout')

wire n774;
// (6, 12, 'lutff_5/lout')

wire n775;
// (6, 4, 'lutff_1/lout')

wire n776;
// (8, 12, 'lutff_7/lout')

wire n777;
// (7, 6, 'lutff_1/lout')

wire n778;
// (9, 6, 'lutff_3/lout')

wire n779;
// (5, 9, 'lutff_4/lout')

wire n780;
// (2, 5, 'lutff_1/out')

wire n781;
// (2, 5, 'lutff_1/lout')

wire n782;
// (6, 5, 'lutff_2/lout')

wire n783;
// (7, 9, 'lutff_6/lout')

wire n784;
// (11, 11, 'lutff_2/lout')

wire n785;
// (8, 5, 'lutff_4/lout')

wire n786;
// (9, 10, 'lutff_0/lout')

wire n787;
// (5, 13, 'lutff_1/lout')

wire n788;
// (7, 10, 'lutff_7/lout')

wire n789;
// (7, 2, 'lutff_3/lout')

wire n790;
// (4, 9, 'lutff_0/lout')

wire n791;
// (8, 9, 'lutff_1/lout')

wire n792;
// (2, 9, 'lutff_7/lout')

wire n793;
// (11, 7, 'lutff_4/lout')

wire n794;
// (4, 6, 'lutff_3/lout')

wire n795;
// (5, 5, 'lutff_2/lout')

wire n796;
// (7, 5, 'lutff_4/lout')

wire n797;
// (6, 12, 'lutff_0/lout')

wire n798;
// (4, 12, 'lutff_1/lout')

wire n799;
// (8, 12, 'lutff_2/lout')

wire n800;
// (6, 4, 'lutff_5/lout')

wire n801;
// (8, 4, 'lutff_7/lout')

wire n802;
// (12, 10, 'lutff_1/lout')

wire n803;
// (7, 6, 'lutff_5/lout')

wire n804;
// (8, 13, 'lutff_3/lout')

wire n805;
// (7, 9, 'lutff_1/lout')

wire n806;
// (9, 9, 'lutff_3/lout')

wire n807;
// (2, 5, 'lutff_5/lout')

wire n808;
// (6, 5, 'lutff_6/lout')

wire n809;
// (7, 10, 'lutff_2/lout')

wire n810;
// (5, 13, 'lutff_5/lout')

wire n811;
// (2, 9, 'lutff_2/lout')

wire n812;
// (7, 2, 'lutff_7/lout')

wire n813;
// (4, 9, 'lutff_4/lout')

wire n814;
// (8, 8, 'lutff_0/lout')

wire n815;
// (6, 8, 'lutff_7/lout')

wire n816;
// (7, 13, 'lutff_3/lout')

wire n817;
// (9, 13, 'lutff_5/lout')

wire n818;
// (5, 5, 'lutff_6/lout')

wire n819;
// (6, 12, 'lutff_4/lout')

wire n820;
// (6, 4, 'lutff_0/lout')

wire n821;
// (8, 12, 'lutff_6/lout')

wire n822;
// (8, 4, 'lutff_2/lout')

wire n823;
// (7, 6, 'lutff_0/lout')

wire n824;
// (5, 9, 'lutff_3/lout')

wire n825;
// (2, 5, 'lutff_0/out')

wire n826;
// (2, 5, 'lutff_0/lout')

wire n827;
// (2, 5, 'carry_in_mux')

// Carry-In for (2 5)
assign n827 = 1;

wire n828;
// (6, 5, 'lutff_1/lout')

wire n829;
// (7, 9, 'lutff_5/lout')

wire n830;
// (8, 5, 'lutff_3/lout')

wire n831;
// (9, 9, 'lutff_7/lout')

wire n832;
// (5, 12, 'lutff_4/lout')

wire n833;
// (6, 8, 'lutff_2/lout')

wire n834;
// (7, 12, 'lutff_6/lout')

wire n835;
// (4, 8, 'lutff_3/lout')

wire n836;
// (8, 8, 'lutff_4/lout')

wire n837;
// (5, 5, 'lutff_1/lout')

wire n838;
// (7, 13, 'lutff_7/lout')

wire n839;
// (7, 5, 'lutff_3/lout')

wire n840;
// (4, 12, 'lutff_0/lout')

wire n841;
// (8, 12, 'lutff_1/lout')

wire n842;
// (6, 4, 'lutff_4/lout')

wire n843;
// (8, 4, 'lutff_6/lout')

wire n844;
// (12, 10, 'lutff_0/lout')

wire n845;
// (6, 7, 'lutff_6/lout')

wire n846;
// (7, 9, 'lutff_0/lout')

wire n847;
// (9, 6, 'lutff_6/lout')

wire n848;
// (1, 6, 'lutff_6/lout')

wire n849;
// (9, 9, 'lutff_2/lout')

wire n850;
// (11, 11, 'lutff_5/lout')

wire n851;
// (1, 3, 'lutff_0/out')

wire n852;
// (1, 3, 'lutff_0/lout')

wire n853;
// (1, 3, 'carry_in_mux')

// Carry-In for (1 3)
assign n853 = 1;

wire n854;
// (6, 11, 'lutff_3/lout')

wire n855;
// (8, 11, 'lutff_5/lout')

wire n856;
// (7, 12, 'lutff_1/lout')

wire n857;
// (9, 12, 'lutff_3/lout')

wire n858;
// (5, 4, 'lutff_4/lout')

wire n859;
// (6, 8, 'lutff_6/lout')

wire n860;
// (7, 4, 'lutff_6/lout')

wire n861;
// (7, 13, 'lutff_2/lout')

wire n862;
// (5, 5, 'lutff_5/lout')

wire n863;
// (7, 5, 'lutff_7/lout')

wire n864;
// (8, 4, 'lutff_1/lout')

wire n865;
// (2, 4, 'lutff_7/lout')

wire n866;
// (6, 7, 'lutff_1/lout')

wire n867;
// (8, 7, 'lutff_3/lout')

wire n868;
// (5, 8, 'lutff_6/lout')

wire n869;
// (9, 8, 'lutff_1/lout')

wire n870;
// (5, 11, 'lutff_2/lout')

wire n871;
// (4, 4, 'lutff_5/lout')

wire n872;
// (7, 11, 'lutff_4/lout')

wire n873;
// (4, 7, 'lutff_1/lout')

wire n874;
// (1, 3, 'lutff_4/lout')

wire n875;
// (8, 11, 'lutff_0/lout')

wire n876;
// (6, 11, 'lutff_7/lout')

wire n877;
// (11, 6, 'lutff_7/lout')

wire n878;
// (11, 9, 'lutff_3/lout')

wire n879;
// (5, 12, 'lutff_3/lout')

wire n880;
// (7, 12, 'lutff_5/lout')

wire n881;
// (6, 8, 'lutff_1/lout')

wire n882;
// (4, 8, 'lutff_2/lout')

wire n883;
// (9, 12, 'lutff_7/lout')

wire n884;
// (8, 8, 'lutff_3/lout')

wire n885;
// (7, 4, 'lutff_1/lout')

wire n886;
// (5, 5, 'lutff_0/lout')

wire n887;
// (7, 5, 'lutff_2/lout')

wire n888;
// (9, 5, 'lutff_4/lout')

wire n889;
// (4, 11, 'lutff_3/lout')

wire n890;
// (2, 3, 'lutff_6/lout')

wire n891;
// (6, 7, 'lutff_5/lout')

wire n892;
// (8, 7, 'lutff_7/lout')

wire n893;
// (5, 8, 'lutff_1/lout')

wire n894;
// (7, 8, 'lutff_3/lout')

wire n895;
// (4, 4, 'lutff_0/lout')

wire n896;
// (9, 8, 'lutff_5/lout')

wire n897;
// (5, 11, 'lutff_6/lout')

wire n898;
// (4, 7, 'lutff_5/lout')

wire n899;
// (6, 11, 'lutff_2/lout')

wire n900;
// (8, 11, 'lutff_4/lout')

wire n901;
// (11, 9, 'lutff_7/lout')

wire n902;
// (7, 12, 'lutff_0/lout')

wire n903;
// (5, 12, 'lutff_7/lout')

wire n904;
// (9, 12, 'lutff_2/lout')

wire n905;
// (7, 4, 'lutff_5/lout')

wire n906;
// (8, 3, 'lutff_5/lout')

wire n907;
// (5, 7, 'lutff_4/lout')

wire n908;
// (2, 3, 'lutff_1/lout')

wire n909;
// (4, 11, 'lutff_7/lout')

wire n910;
// (7, 7, 'lutff_6/lout')

wire n911;
// (4, 14, 'lutff_3/lout')

wire n912;
// (8, 7, 'lutff_2/lout')

wire n913;
// (11, 5, 'lutff_5/lout')

wire n914;
// (5, 8, 'lutff_5/lout')

wire n915;
// (9, 8, 'lutff_0/lout')

wire n916;
// (7, 8, 'lutff_7/lout')

wire n917;
// (5, 11, 'lutff_1/lout')

wire n918;
// (4, 4, 'lutff_4/lout')

wire n919;
// (7, 11, 'lutff_3/lout')

wire n920;
// (4, 7, 'lutff_0/lout')

wire n921;
// (1, 3, 'lutff_3/lout')

wire n922;
// (2, 7, 'lutff_7/lout')

wire n923;
// (11, 9, 'lutff_2/lout')

wire n924;
// (5, 12, 'lutff_2/lout')

wire n925;
// (4, 8, 'lutff_1/lout')

wire n926;
// (9, 12, 'lutff_6/lout')

wire n927;
// (7, 4, 'lutff_0/lout')

wire n928;
// (2, 11, 'lutff_4/lout')

wire n929;
// (12, 11, 'lutff_7/lout')

wire n930;
// (8, 3, 'lutff_0/lout')

wire n931;
// (6, 3, 'lutff_7/lout')

wire n932;
// (4, 11, 'lutff_2/lout')

wire n933;
// (7, 7, 'lutff_1/lout')

wire n934;
// (2, 3, 'lutff_5/lout')

wire n935;
// (6, 7, 'lutff_4/lout')

wire n936;
// (8, 7, 'lutff_6/lout')

wire n937;
// (5, 8, 'lutff_0/lout')

wire n938;
// (7, 8, 'lutff_2/lout')

wire n939;
// (12, 12, 'lutff_7/lout')

wire n940;
// (9, 8, 'lutff_4/lout')

wire n941;
// (5, 11, 'lutff_5/lout')

wire n942;
// (7, 11, 'lutff_7/lout')

wire n943;
// (4, 7, 'lutff_4/lout')

wire n944;
// (11, 6, 'lutff_1/lout')

wire n945;
// (5, 14, 'lutff_7/lout')

wire n946;
// (6, 10, 'lutff_5/lout')

wire n947;
// (11, 9, 'lutff_6/lout')

wire n948;
// (8, 10, 'lutff_7/lout')

wire n949;
// (6, 13, 'lutff_1/lout')

wire n950;
// (8, 2, 'lutff_3/lout')

wire n951;
// (9, 11, 'lutff_5/lout')

wire n952;
// (12, 11, 'lutff_2/lout')

wire n953;
// (5, 6, 'lutff_2/lout')

wire n954;
// (4, 10, 'lutff_5/lout')

wire n955;
// (6, 3, 'lutff_2/lout')

wire n956;
// (8, 3, 'lutff_4/lout')

wire n957;
// (11, 12, 'lutff_7/lout')

wire n958;
// (2, 3, 'lutff_0/lout')

wire n959;
// (7, 7, 'lutff_5/lout')

wire n960;
// (4, 3, 'lutff_2/lout')

wire n961;
// (8, 7, 'lutff_1/lout')

wire n962;
// (11, 5, 'lutff_4/lout')

wire n963;
// (8, 6, 'lutff_5/lout')

wire n964;
// (5, 11, 'lutff_0/lout')

wire n965;
// (7, 11, 'lutff_2/lout')

wire n966;
// (2, 6, 'lutff_1/lout')

wire n967;
// (5, 14, 'lutff_2/lout')

wire n968;
// (6, 10, 'lutff_0/lout')

wire n969;
// (7, 14, 'lutff_4/lout')

wire n970;
// (11, 9, 'lutff_1/lout')

wire n971;
// (8, 10, 'lutff_2/lout')

wire n972;
// (9, 14, 'lutff_6/lout')

wire n973;
// (6, 13, 'lutff_5/lout')

wire n974;
// (8, 2, 'lutff_7/lout')

wire n975;
// (7, 3, 'lutff_3/lout')

wire n976;
// (4, 10, 'lutff_0/lout')

wire n977;
// (2, 10, 'lutff_7/lout')

wire n978;
// (5, 6, 'lutff_6/lout')

wire n979;
// (6, 14, 'lutff_6/lout')

wire n980;
// (6, 3, 'lutff_6/lout')

wire n981;
// (4, 2, 'lutff_5/lout')

wire n982;
// (6, 6, 'lutff_2/lout')

wire n983;
// (7, 15, 'lutff_4/lout')

wire n984;
// (4, 11, 'lutff_1/lout')

wire n985;
// (7, 7, 'lutff_0/lout')

wire n986;
// (2, 3, 'lutff_4/lout')

wire n987;
// (8, 6, 'lutff_0/lout')

wire n988;
// (6, 9, 'lutff_3/lout')

wire n989;
// (8, 9, 'lutff_5/lout')

wire n990;
// (2, 6, 'lutff_5/lout')

wire n991;
// (5, 14, 'lutff_6/lout')

wire n992;
// (9, 14, 'lutff_1/lout')

wire n993;
// (4, 6, 'lutff_7/lout')

wire n994;
// (6, 10, 'lutff_4/lout')

wire n995;
// (8, 10, 'lutff_6/lout')

wire n996;
// (6, 13, 'lutff_0/lout')

wire n997;
// (11, 8, 'lutff_0/lout')

wire n998;
// (8, 2, 'lutff_2/lout')

wire n999;
// (2, 10, 'lutff_2/lout')

wire n1000;
// (7, 3, 'lutff_7/lout')

wire n1001;
// (4, 10, 'lutff_4/lout')

wire n1002;
// (8, 14, 'lutff_3/lout')

wire n1003;
// (11, 12, 'lutff_6/lout')

wire n1004;
// (8, 13, 'lutff_7/lout')

wire n1005;
// (7, 7, 'lutff_4/lout')

wire n1006;
// (5, 10, 'lutff_4/lout')

wire n1007;
// (5, 13, 'lutff_0/lout')

wire n1008;
// (7, 10, 'lutff_6/lout')

wire n1009;
// (8, 6, 'lutff_4/lout')

wire n1010;
// (7, 2, 'lutff_2/lout')

wire n1011;
// (8, 9, 'lutff_0/lout')

wire n1012;
// (1, 5, 'lutff_2/lout')

wire n1013;
// (6, 9, 'lutff_7/lout')

wire n1014;
// (2, 6, 'lutff_0/lout')

wire n1015;
// (5, 14, 'lutff_1/lout')

wire n1016;
// (4, 6, 'lutff_2/lout')

wire n1017;
// (7, 14, 'lutff_3/lout')

wire n1018;
// (8, 10, 'lutff_1/lout')

wire n1019;
// (9, 14, 'lutff_5/lout')

wire n1020;
// (6, 13, 'lutff_4/lout')

wire n1021;
// (8, 2, 'lutff_6/lout')

wire n1022;
// (11, 8, 'lutff_4/lout')

wire n1023;
// (7, 3, 'lutff_2/lout')

wire n1024;
// (2, 10, 'lutff_6/lout')

wire n1025;
// (5, 6, 'lutff_5/lout')

wire n1026;
// (12, 11, 'lutff_5/lout')

wire n1027;
// (2, 2, 'lutff_2/lout')

wire n1028;
// (7, 6, 'lutff_4/lout')

wire n1029;
// (11, 12, 'lutff_1/lout')

wire n1030;
// (8, 13, 'lutff_2/lout')

wire n1031;
// (5, 9, 'lutff_7/lout')

wire n1032;
// (2, 5, 'lutff_4/lout')

wire n1033;
// (6, 5, 'lutff_5/lout')

wire n1034;
// (8, 5, 'lutff_7/lout')

wire n1035;
// (7, 10, 'lutff_1/lout')

wire n1036;
// (5, 13, 'lutff_4/lout')

wire n1037;
// (6, 9, 'lutff_2/lout')

wire n1038;
// (7, 2, 'lutff_6/lout')

wire n1039;
// (4, 9, 'lutff_3/lout')

wire n1040;
// (8, 9, 'lutff_4/lout')

wire n1041;
// (11, 7, 'lutff_7/lout')

wire n1042;
// (4, 6, 'lutff_6/lout')

wire n1043;
// (8, 2, 'lutff_1/lout')

wire n1044;
// (6, 12, 'lutff_3/lout')

wire n1045;
// (8, 12, 'lutff_5/lout')

wire n1046;
// (5, 6, 'lutff_0/lout')

wire n1047;
// (5, 9, 'lutff_2/lout')

wire n1048;
// (6, 5, 'lutff_0/lout')

wire n1049;
// (8, 13, 'lutff_6/lout')

wire n1050;
// (4, 5, 'lutff_1/lout')

wire n1051;
// (9, 9, 'lutff_6/lout')

wire n1052;
// (7, 9, 'lutff_4/lout')

wire n1053;
// (8, 5, 'lutff_2/lout')

wire n1054;
// (11, 3, 'lutff_5/lout')

wire n1055;
// (5, 10, 'lutff_3/lout')

wire n1056;
// (7, 10, 'lutff_5/lout')

wire n1057;
// (8, 6, 'lutff_3/lout')

wire n1058;
// (7, 2, 'lutff_1/lout')

wire n1059;
// (6, 9, 'lutff_6/lout')

wire n1060;
// (4, 9, 'lutff_7/lout')

wire n1061;
// (11, 7, 'lutff_2/lout')

wire n1062;
// (5, 14, 'lutff_0/lout')

wire n1063;
// (4, 6, 'lutff_1/lout')

wire n1064;
// (7, 14, 'lutff_2/lout')

wire n1065;
// (9, 14, 'lutff_4/lout')

wire n1066;
// (7, 13, 'lutff_6/lout')

wire n1067;
// (11, 8, 'lutff_3/lout')

wire n1068;
// (8, 12, 'lutff_0/lout')

wire n1069;
// (6, 12, 'lutff_7/lout')

wire n1070;
// (6, 4, 'lutff_3/lout')

wire n1071;
// (8, 4, 'lutff_5/lout')

wire n1072;
// (7, 6, 'lutff_3/lout')

wire n1073;
// (8, 13, 'lutff_1/lout')

wire n1074;
// (5, 9, 'lutff_6/lout')

wire n1075;
// (9, 9, 'lutff_1/lout')

wire n1076;
// (2, 5, 'lutff_3/lout')

wire n1077;
// (6, 5, 'lutff_4/lout')

wire n1078;
// (11, 11, 'lutff_4/lout')

wire n1079;
// (8, 5, 'lutff_6/lout')

wire n1080;
// (7, 10, 'lutff_0/lout')

wire n1081;
// (5, 10, 'lutff_7/lout')

wire n1082;
// (5, 13, 'lutff_3/lout')

wire n1083;
// (2, 9, 'lutff_0/lout')

wire n1084;
// (7, 2, 'lutff_5/lout')

wire n1085;
// (4, 9, 'lutff_2/lout')

wire n1086;
// (8, 9, 'lutff_3/lout')

wire n1087;
// (6, 8, 'lutff_5/lout')

wire n1088;
// (8, 8, 'lutff_7/lout')

wire n1089;
// (9, 13, 'lutff_3/lout')

wire n1090;
// (5, 5, 'lutff_4/lout')

wire n1091;
// (6, 12, 'lutff_2/lout')

wire n1092;
// (7, 5, 'lutff_6/lout')

wire n1093;
// (8, 12, 'lutff_4/lout')

wire n1094;
// (8, 4, 'lutff_0/lout')

wire n1095;
// (6, 4, 'lutff_7/lout')

wire n1096;
// (7, 6, 'lutff_7/lout')

wire n1097;
// (5, 9, 'lutff_1/lout')

wire n1098;
// (7, 9, 'lutff_3/lout')

wire n1099;
// (4, 5, 'lutff_0/lout')

wire n1100;
// (9, 9, 'lutff_5/lout')

wire n1101;
// (2, 5, 'lutff_7/lout')

wire n1102;
// (8, 5, 'lutff_1/lout')

wire n1103;
// (7, 2, 'lutff_0/lout')

wire n1104;
// (11, 7, 'lutff_1/lout')

wire n1105;
// (8, 8, 'lutff_2/lout')

wire n1106;
// (7, 13, 'lutff_5/lout')

wire n1107;
// (7, 5, 'lutff_1/lout')

wire n1108;
// (9, 13, 'lutff_7/lout')

wire n1109;
// (6, 12, 'lutff_6/lout')

wire n1110;
// (6, 4, 'lutff_2/lout')

wire n1111;
// (8, 4, 'lutff_4/lout')

wire n1112;
// (7, 6, 'lutff_2/lout')

wire n1113;
// (9, 9, 'lutff_0/lout')

wire n1114;
// (2, 5, 'lutff_2/lout')

wire n1115;
// (11, 11, 'lutff_3/lout')

wire n1116;
// (6, 11, 'lutff_1/lout')

wire n1117;
// (8, 11, 'lutff_3/lout')

assign n627  = /* LUT    1  3  1 */ 1'b0;
assign n781  = /* LUT    2  5  1 */ 1'b0;
assign n826  = /* LUT    2  5  0 */ 1'b0;
assign n852  = /* LUT    1  3  0 */ 1'b0;
assign n561  = /* LUT    5 12  6 */ n213;
assign n562  = /* LUT    9 12  1 */ (n471 ? (n31 ? n517 : 1'b0) : (n31 ? !n517 : 1'b1));
assign n563  = /* LUT    2  8  3 */ !rst;
assign n564  = /* LUT    6  8  4 */ (n192 ? (n122 ? 1'b1 : !n260) : (n122 ? (n288 ? !n260 : n260) : !n288));
assign n565  = /* LUT    4  8  5 */ n123;
assign n566  = /* LUT    8  8  6 */ (n30 ? (n443 ? n441 : !n441) : (n443 ? !n441 : n441));
assign n567  = /* LUT    7  4  4 */ (n158 ? !n236 : n236);
assign n568  = /* LUT    1  7  4 */ n72;
assign n569  = /* LUT    7 13  0 */ (n286 ? n395 : (n340 ? n372 : !n372));
assign n570  = /* LUT    9 13  2 */ n530;
assign n571  = /* LUT    5  5  3 */ (n154 ? 1'b0 : !n157);
assign n572  = /* LUT    7  5  5 */ (n170 ? (n21 ? 1'b0 : (n19 ? !n22 : 1'b1)) : 1'b0);
assign n573  = /* LUT    4 12  2 */ n208;
assign n574  = /* LUT    8 12  3 */ n472;
assign n575  = /* LUT    9  5  7 */ n531;
assign n576  = /* LUT    6  4  6 */ (n230 ? 1'b0 : !n234);
assign n577  = /* LUT    5  9  0 */ n191;
assign n578  = /* LUT    7  9  2 */ (n35 ? (n96 ? n88 : 1'b1) : (n96 ? !n88 : 1'b0));
assign n579  = /* LUT    9  9  4 */ (n445 ? (n31 ? n498 : 1'b0) : (n31 ? !n498 : 1'b1));
assign n580  = /* LUT    5  8  4 */ n174;
assign n581  = /* LUT    7  8  6 */ (n339 ? (n255 ? (n346 ? 1'b1 : n193) : (n346 ? n193 : 1'b1)) : (n255 ? 1'b0 : n193));
assign n582  = /* LUT    1  3  2 */ (n57 ? (n6 ? 1'b0 : !n51) : (n6 ? !n51 : 1'b0));
assign n583  = /* LUT    8 11  7 */ (n25 ? (n68 ? n477 : n464) : n477);
assign n584  = /* LUT   11  6  5 */ n535;
assign n585  = /* LUT    5 12  1 */ n168;
assign n586  = /* LUT    7 12  3 */ n42;
assign n587  = /* LUT    9 12  5 */ (n70 ? n485 : n532);
assign n588  = /* LUT    8  8  1 */ (n349 ? !n425 : n425);
assign n589  = /* LUT    7 13  4 */ n385;
assign n590  = /* LUT    7  5  0 */ (n330 ? (n21 ? (n22 ? 1'b0 : !n63) : n22) : 1'b0);
assign n591  = /* LUT    9 13  6 */ n522;
assign n592  = /* LUT    5  5  7 */ n148;
assign n593  = /* LUT    9  5  2 */ n489;
assign n594  = /* LUT   12  9  5 */ n546;
assign n595  = /* LUT    4 12  6 */ n143;
assign n596  = /* LUT    8  4  3 */ (n414 ? (n416 ? !n171 : n171) : (n416 ? n171 : !n171));
assign n597  = /* LUT    6  7  3 */ (n266 ? (n254 ? (n261 ? n192 : !n192) : (n261 ? !n192 : n192)) : (n254 ? (n261 ? !n192 : n192) : (n261 ? n192 : !n192)));
assign n598  = /* LUT    8  7  5 */ (n433 ? (n431 ? (n254 ? !n429 : 1'b1) : (n254 ? n429 : 1'b0)) : (n431 ? (n254 ? n429 : 1'b0) : (n254 ? !n429 : 1'b1)));
assign n599  = /* LUT    7  8  1 */ (n262 ? (n352 ? !n261 : 1'b1) : (n352 ? (n261 ? !n348 : n348) : !n348));
assign n600  = /* LUT    9  8  3 */ (n496 ? (n493 ? (n418 ? 1'b1 : n88) : (n418 ? n88 : 1'b1)) : (n493 ? (n418 ? 1'b0 : !n88) : (n418 ? !n88 : 1'b0)));
assign n601  = /* LUT    5 11  4 */ n203;
assign n602  = /* LUT    7 11  6 */ n368;
assign n603  = /* LUT    4  7  3 */ n117;
assign n604  = /* LUT    6 11  0 */ (n293 ? (n107 ? (n360 ? !n286 : 1'b1) : (n360 ? 1'b1 : !n286)) : 1'b0);
assign n605  = /* LUT   11  6  0 */ (select ? !n538 : 1'b0);
assign n606  = /* LUT    8 11  2 */ (n176 ? (n31 ? n454 : 1'b0) : (n31 ? !n454 : 1'b1));
assign n607  = /* LUT   11  9  5 */ (n440 ? (n31 ? !n549 : 1'b1) : (n31 ? n549 : 1'b0));
assign n608  = /* LUT    9 12  0 */ (n70 ? !n517 : !n514);
assign n609  = /* LUT    6  8  3 */ (n122 ? (n276 ? (n287 ? n196 : !n196) : (n287 ? !n196 : n196)) : (n276 ? (n287 ? !n196 : n196) : (n287 ? n196 : !n196)));
assign n610  = /* LUT    7 12  7 */ n377;
assign n611  = /* LUT    4  8  4 */ n126;
assign n612  = /* LUT    7  4  3 */ (n158 ? (n329 ? !n155 : n155) : (n329 ? n155 : !n155));
assign n613  = /* LUT    8  8  5 */ (n350 ? (n431 ? (n427 ? n436 : !n436) : (n427 ? !n436 : n436)) : (n431 ? (n427 ? !n436 : n436) : (n427 ? n436 : !n436)));
assign n614  = /* LUT   11 10  6 */ n518;
assign n615  = /* LUT    8  3  3 */ (n322 ? (n404 ? n324 : 1'b1) : (n404 ? (n324 ? n400 : !n400) : !n400));
assign n616  = /* LUT    6  6  6 */ n340;
assign n617  = /* LUT    8  7  0 */ (n426 ? (n254 ? !n27 : n27) : 1'b0);
assign n618  = /* LUT    6  7  7 */ (n254 ? n261 : !n261);
assign n619  = /* LUT   11 13  7 */ n383;
assign n620  = /* LUT   11  5  3 */ n536;
assign n621  = /* LUT    1  6  7 */ n23;
assign n622  = /* LUT    5  8  3 */ n180;
assign n623  = /* LUT    7  8  5 */ (n261 ? (n276 ? (n254 ? 1'b0 : !n260) : (n254 ? 1'b1 : n260)) : (n254 ? !n260 : 1'b0));
assign n624  = /* LUT    7 11  1 */ (n367 ? (n167 ? (n470 ? !n286 : 1'b1) : (n470 ? 1'b1 : !n286)) : 1'b0);
assign n625  = /* LUT    9  8  7 */ n492;
assign n628  = /* LUT    6 11  4 */ (n286 ? n43 : (n107 ? n360 : !n360));
assign n629  = /* LUT   11  6  4 */ n417;
assign n630  = /* LUT    8 11  6 */ (n70 ? n454 : n146);
assign n631  = /* LUT   11  9  0 */ (select ? 1'b1 : n547);
assign n632  = /* LUT    5 12  0 */ n167;
assign n633  = /* LUT    7 12  2 */ (n25 ? (n68 ? n371 : n365) : n371);
assign n634  = /* LUT    9 12  4 */ (n70 ? n87 : n513);
assign n635  = /* LUT    5  4  5 */ n101;
assign n636  = /* LUT    7  4  7 */ (n233 ? !n322 : n322);
assign n637  = /* LUT   11 10  1 */ (select ? 1'b1 : n458);
assign n638  = /* LUT    6  6  1 */ n107;
assign n639  = /* LUT    8  3  7 */ (n325 ? (n235 ? 1'b1 : n249) : (n235 ? (n403 ? n249 : !n249) : n403));
assign n640  = /* LUT    4 11  0 */ n141;
assign n641  = /* LUT    2  3  3 */ (n1 ? (n9 ? 1'b1 : rst) : 1'b1);
assign n642  = /* LUT    2 14  3 */ n47;
assign n643  = /* LUT    4  3  5 */ (rst ? 1'b0 : (n4 ? 1'b1 : (n60 ? !n12 : 1'b0)));
assign n644  = /* LUT    6  7  2 */ (n263 ? (n258 ? (n256 ? n257 : 1'b1) : (n256 ? !n257 : 1'b0)) : (n258 ? (n256 ? !n257 : 1'b0) : (n256 ? n257 : 1'b1)));
assign n645  = /* LUT    8  7  4 */ (n276 ? (n426 ? !n347 : 1'b0) : (n426 ? (n347 ? !n429 : n429) : n429));
assign n646  = /* LUT    7  8  0 */ (n346 ? (n339 ? (n193 ? 1'b0 : n255) : n193) : (n339 ? (n193 ? 1'b0 : !n255) : 1'b1));
assign n647  = /* LUT    5  8  7 */ n124;
assign n648  = /* LUT    9  8  2 */ n509;
assign n649  = /* LUT    5 11  3 */ n205;
assign n650  = /* LUT    7 11  5 */ n364;
assign n651  = /* LUT    4  7  2 */ n120;
assign n652  = /* LUT    8 11  1 */ n467;
assign n653  = /* LUT    6 10  3 */ n281;
assign n654  = /* LUT   11  9  4 */ (n440 ? (n137 ? (n546 ? n31 : 1'b0) : (n546 ? !n31 : 1'b1)) : (n137 ? (n546 ? !n31 : 1'b1) : (n546 ? n31 : 1'b0)));
assign n655  = /* LUT    8 10  5 */ (n446 ? !n72 : n72);
assign n656  = /* LUT    5  4  0 */ (n151 ? (n10 ? 1'b1 : (n11 ? 1'b1 : n49)) : 1'b0);
assign n657  = /* LUT    7  4  2 */ (n155 ? !n236 : n236);
assign n658  = /* LUT    9 11  3 */ n508;
assign n659  = /* LUT    2 10  1 */ n80;
assign n660  = /* LUT    7  3  6 */ (n320 ? (n318 ? (n325 ? 1'b1 : n248) : (n325 ? 1'b0 : !n248)) : (n318 ? (n325 ? 1'b0 : !n248) : (n325 ? 1'b1 : n248)));
assign n661  = /* LUT    6  3  0 */ (n149 ? 1'b0 : !n229);
assign n662  = /* LUT    8  3  2 */ (n324 ? (n404 ? n322 : 1'b1) : (n404 ? (n322 ? !n402 : n402) : n402));
assign n663  = /* LUT    2  2  6 */ (rst ? 1'b1 : (n9 ? !n52 : 1'b0));
assign n664  = /* LUT    6  6  5 */ n168;
assign n665  = /* LUT    9  4  0 */ n14;
assign n666  = /* LUT    7 15  7 */ n390;
assign n667  = /* LUT    4 11  4 */ n142;
assign n668  = /* LUT    7  7  3 */ (n257 ? (n256 ? (n183 ? !n184 : 1'b0) : (n183 ? 1'b0 : !n184)) : (n256 ? (n183 ? n184 : 1'b0) : (n183 ? 1'b0 : n184)));
assign n669  = /* LUT    4  3  0 */ (n60 ? 1'b0 : (n10 ? 1'b0 : (n11 ? 1'b0 : !n4)));
assign n670  = /* LUT    9  7  5 */ n501;
assign n671  = /* LUT    2  3  7 */ (n56 ? 1'b0 : (n59 ? (n9 ? 1'b1 : n60) : 1'b1));
assign n672  = /* LUT    5  8  2 */ n181;
assign n673  = /* LUT    7  8  4 */ (n260 ? (n352 ? n192 : 1'b0) : (n352 ? (n351 ? !n192 : n192) : !n351));
assign n674  = /* LUT    7 11  0 */ (n70 ? !n369 : !n379);
assign n675  = /* LUT    5 11  7 */ (n25 ? (n68 ? n85 : n194) : n85);
assign n676  = /* LUT    8 10  0 */ (n28 ? (n31 ? !n455 : 1'b1) : (n31 ? n455 : 1'b0));
assign n677  = /* LUT    6 10  7 */ n101;
assign n678  = /* LUT    6 13  3 */ n301;
assign n679  = /* LUT    8  2  5 */ (n398 ? (n306 ? (n312 ? n308 : !n308) : (n312 ? 1'b0 : n308)) : (n306 ? (n312 ? !n308 : 1'b0) : 1'b1));
assign n680  = /* LUT    9 11  7 */ (n528 ? (n518 ? n88 : 1'b1) : (n518 ? !n88 : 1'b0));
assign n681  = /* LUT    7  3  1 */ (n319 ? n318 : !n318);
assign n682  = /* LUT    9  3  3 */ n487;
assign n683  = /* LUT    5  6  4 */ n166;
assign n684  = /* LUT    2  2  1 */ (n49 ? !n55 : 1'b0);
assign n685  = /* LUT    6  3  4 */ (n231 ? (n10 ? 1'b1 : (n11 ? 1'b1 : n49)) : 1'b0);
assign n686  = /* LUT    4 10  7 */ (n130 ? (n72 ? n88 : 1'b1) : (n72 ? !n88 : 1'b0));
assign n687  = /* LUT    8  3  6 */ (n305 ? (n410 ? (n399 ? n152 : 1'b1) : (n399 ? !n152 : 1'b0)) : (n410 ? (n399 ? !n152 : 1'b0) : (n399 ? n152 : 1'b1)));
assign n688  = /* LUT   11 12  0 */ (n471 ? (n516 ? n31 : 1'b0) : (n516 ? !n31 : 1'b1));
assign n689  = /* LUT    7 15  2 */ n396;
assign n690  = /* LUT   11  4  5 */ n115;
assign n691  = /* LUT    5  7  5 */ n71;
assign n692  = /* LUT    2  3  2 */ (n56 ? (n8 ? (n7 ? n6 : 1'b0) : 1'b0) : 1'b0);
assign n693  = /* LUT    7  7  7 */ (n343 ? (n344 ? n342 : !n342) : (n344 ? !n342 : n342));
assign n694  = /* LUT    8  6  7 */ (n257 ? (n184 ? 1'b1 : n430) : (n184 ? n428 : (n430 ? n428 : !n428)));
assign n695  = /* LUT    6  9  1 */ (n265 ? n359 : !n359);
assign n696  = /* LUT    2  6  3 */ (n19 ? (n22 ? (n63 ? 1'b0 : !n21) : 1'b0) : 1'b0);
assign n697  = /* LUT    5 14  4 */ (n25 ? (n68 ? n222 : n221) : n222);
assign n698  = /* LUT    6 10  2 */ n282;
assign n699  = /* LUT    7 14  6 */ n393;
assign n700  = /* LUT    8 10  4 */ (n70 ? n460 : n505);
assign n701  = /* LUT    8  2  0 */ (n310 ? n406 : !n406);
assign n702  = /* LUT    6 13  7 */ (n25 ? (n68 ? n298 : n296) : n298);
assign n703  = /* LUT    6  2  7 */ (n227 ? n152 : !n152);
assign n704  = /* LUT   11  8  7 */ n552;
assign n705  = /* LUT    9 11  2 */ n507;
assign n706  = /* LUT    2 10  0 */ n79;
assign n707  = /* LUT    7  3  5 */ (n233 ? n326 : !n326);
assign n708  = /* LUT    4 10  2 */ n136;
assign n709  = /* LUT    9  3  7 */ n238;
assign n710  = /* LUT    8  3  1 */ (n235 ? (n325 ? 1'b0 : (n314 ? n248 : !n248)) : (n325 ? (n314 ? n248 : !n248) : 1'b0));
assign n711  = /* LUT    4  2  7 */ (rst ? 1'b0 : !n103);
assign n712  = /* LUT    7  7  2 */ (n342 ? (n341 ? (n257 ? !n256 : 1'b0) : (n257 ? n256 : 1'b1)) : (n341 ? (n257 ? n256 : 1'b1) : (n257 ? !n256 : 1'b0)));
assign n713  = /* LUT    5 10  2 */ (n195 ? (n148 ? (n38 ? !n286 : 1'b1) : (n38 ? 1'b1 : !n286)) : 1'b0);
assign n714  = /* LUT    7 10  4 */ (n361 ? (n228 ? (n462 ? !n286 : 1'b1) : (n462 ? 1'b1 : !n286)) : 1'b0);
assign n715  = /* LUT   11  5  1 */ (n534 ? (n115 ? n88 : 1'b1) : (n115 ? !n88 : 1'b0));
assign n716  = /* LUT    8  6  2 */ (n346 ? (n255 ? 1'b0 : !n339) : (n255 ? 1'b1 : n193));
assign n717  = /* LUT    6  9  5 */ (n359 ? (n288 ? !n196 : n196) : (n288 ? n196 : !n196));
assign n718  = /* LUT    4  9  6 */ n128;
assign n719  = /* LUT    8  9  7 */ (n70 ? n447 : n504);
assign n720  = /* LUT    4  6  0 */ (n4 ? (n63 ? (n19 ? n109 : 1'b0) : 1'b0) : 1'b0);
assign n721  = /* LUT    7 14  1 */ (n388 ? (n25 ? (n68 ? !n395 : 1'b1) : 1'b1) : 1'b0);
assign n722  = /* LUT    2  6  7 */ (n13 ? 1'b1 : (n61 ? (n20 ? 1'b1 : n62) : 1'b0));
assign n723  = /* LUT    9 14  3 */ n529;
assign n724  = /* LUT    6 10  6 */ n278;
assign n725  = /* LUT    6  2  2 */ (n88 ? !n49 : 1'b0);
assign n726  = /* LUT    6 13  2 */ n297;
assign n727  = /* LUT   11  8  2 */ (n273 ? n115 : !n115);
assign n728  = /* LUT    8  2  4 */ (n308 ? (n312 ? (n306 ? 1'b1 : n398) : (n306 ? n398 : 1'b1)) : (n312 ? 1'b0 : n398));
assign n729  = /* LUT    7  3  0 */ (n227 ? (n325 ? !n248 : 1'b1) : (n326 ? (n325 ? !n248 : 1'b1) : (n325 ? n248 : 1'b0)));
assign n730  = /* LUT    9 11  6 */ (n440 ? !n518 : n518);
assign n731  = /* LUT    2 10  4 */ n77;
assign n732  = /* LUT    5  6  3 */ (n176 ? n163 : !n163);
assign n733  = /* LUT    4 10  6 */ n133;
assign n734  = /* LUT    8 13  0 */ (n70 ? !n483 : !n480);
assign n735  = /* LUT    6  5  3 */ (n10 ? 1'b0 : (n11 ? 1'b0 : !n49));
assign n736  = /* LUT    8  5  5 */ (n169 ? (n253 ? !n408 : n408) : (n253 ? n408 : !n408));
assign n737  = /* LUT    5 10  6 */ n199;
assign n738  = /* LUT    9 10  1 */ n451;
assign n739  = /* LUT    5 13  2 */ (n216 ? (n25 ? (n68 ? !n221 : 1'b1) : 1'b1) : 1'b0);
assign n740  = /* LUT    6  9  0 */ (n265 ? (n122 ? n276 : !n276) : (n122 ? !n276 : n276));
assign n741  = /* LUT    8  6  6 */ (n193 ? (n346 ? (n255 ? n339 : !n339) : n255) : (n346 ? n339 : (n255 ? n339 : !n339)));
assign n742  = /* LUT    4  9  1 */ n24;
assign n743  = /* LUT    8  9  2 */ (n176 ? (n444 ? (n451 ? n31 : 1'b0) : (n451 ? !n31 : 1'b1)) : (n444 ? (n451 ? !n31 : 1'b1) : (n451 ? n31 : 1'b0)));
assign n744  = /* LUT    7  2  4 */ (n318 ? (n304 ? !n316 : n316) : (n304 ? n316 : !n316));
assign n745  = /* LUT   11  7  5 */ n539;
assign n746  = /* LUT    2  6  2 */ (rst ? 1'b1 : (n66 ? 1'b1 : n52));
assign n747  = /* LUT    4  6  4 */ (n4 ? (n109 ? (n19 ? !n63 : 1'b0) : 1'b0) : 1'b0);
assign n748  = /* LUT    7 14  5 */ (n68 ? (n25 ? n386 : n395) : n386);
assign n749  = /* LUT    6 10  1 */ n363;
assign n750  = /* LUT    8 10  3 */ (n70 ? n455 : n457);
assign n751  = /* LUT    6 13  6 */ (n68 ? (n25 ? n218 : n296) : n218);
assign n752  = /* LUT    9 11  1 */ n510;
assign n753  = /* LUT    7  3  4 */ (n315 ? (n160 ? (n161 ? !n324 : n324) : !n324) : (n160 ? 1'b1 : !n161));
assign n754  = /* LUT    4 10  1 */ n135;
assign n755  = /* LUT    5  6  7 */ n165;
assign n756  = /* LUT    2  2  4 */ (rst ? 1'b0 : (n11 ? 1'b1 : (n10 ? !n50 : 1'b0)));
assign n757  = /* LUT    7  6  6 */ (n4 ? (n335 ? (n22 ? !n21 : n21) : 1'b0) : 1'b0);
assign n758  = /* LUT   11 12  3 */ (n273 ? (n31 ? n485 : 1'b0) : (n31 ? !n485 : 1'b1));
assign n759  = /* LUT    8 13  4 */ (n446 ? (n275 ? (n481 ? n31 : 1'b0) : (n481 ? !n31 : 1'b1)) : (n275 ? (n481 ? !n31 : 1'b1) : (n481 ? n31 : 1'b0)));
assign n760  = /* LUT    8  5  0 */ (n59 ? (n420 ? (n412 ? !n423 : n423) : (n412 ? n423 : !n423)) : 1'b0);
assign n761  = /* LUT    2  5  6 */ (n93 ? !n21 : n21);
assign n762  = /* LUT    6  5  7 */ (n232 ? (n242 ? 1'b1 : n241) : (n242 ? 1'b0 : !n241));
assign n763  = /* LUT    5 10  1 */ (n200 ? (n25 ? (n68 ? !n194 : 1'b1) : 1'b1) : 1'b0);
assign n764  = /* LUT    7 10  3 */ (n25 ? (n68 ? 1'b1 : !n371) : (n68 ? !n277 : 1'b1));
assign n765  = /* LUT    8  6  1 */ (n257 ? (n184 ? 1'b0 : !n428) : (n184 ? (n430 ? !n428 : n428) : !n430));
assign n766  = /* LUT    2  9  3 */ n84;
assign n767  = /* LUT    6  9  4 */ (n267 ? (n25 ? (n68 ? !n98 : 1'b1) : 1'b1) : 1'b0);
assign n768  = /* LUT    4  9  5 */ n148;
assign n769  = /* LUT    8  9  6 */ (n176 ? (n440 ? (n31 ? !n448 : 1'b1) : (n31 ? n448 : 1'b0)) : (n440 ? (n31 ? n448 : 1'b0) : (n31 ? !n448 : 1'b1)));
assign n770  = /* LUT   11  7  0 */ n358;
assign n771  = /* LUT    7 14  0 */ (n25 ? (n68 ? 1'b1 : !n392) : (n68 ? !n386 : 1'b1));
assign n772  = /* LUT    2  6  6 */ (n13 ? (n20 ? 1'b1 : n62) : (n20 ? n62 : 1'b1));
assign n773  = /* LUT   11  8  1 */ (select ? 1'b1 : n544);
assign n774  = /* LUT    6 12  5 */ (n286 ? n296 : (n168 ? n366 : !n366));
assign n775  = /* LUT    6  4  1 */ (n149 ? (n230 ? 1'b1 : n234) : (n230 ? n229 : (n234 ? n229 : !n229)));
assign n776  = /* LUT    8 12  7 */ n474;
assign n777  = /* LUT    7  6  1 */ (n32 ? !n331 : n331);
assign n778  = /* LUT    9  6  3 */ n96;
assign n779  = /* LUT    5  9  4 */ n33;
assign n782  = /* LUT    6  5  2 */ (n240 ? (n10 ? 1'b1 : (n11 ? 1'b1 : n49)) : 1'b0);
assign n783  = /* LUT    7  9  6 */ n356;
assign n784  = /* LUT   11 11  2 */ (select ? 1'b1 : n478);
assign n785  = /* LUT    8  5  4 */ (n59 ? (n171 ? (n419 ? n175 : !n175) : (n419 ? !n175 : n175)) : 1'b0);
assign n786  = /* LUT    9 10  0 */ n459;
assign n787  = /* LUT    5 13  1 */ (n25 ? (n68 ? 1'b1 : !n222) : (n68 ? !n220 : 1'b1));
assign n788  = /* LUT    7 10  7 */ (n68 ? (n25 ? n277 : n365) : n277);
assign n789  = /* LUT    7  2  3 */ (n321 ? (n309 ? 1'b0 : (n306 ? n311 : 1'b1)) : 1'b0);
assign n790  = /* LUT    4  9  0 */ n129;
assign n791  = /* LUT    8  9  1 */ (n437 ? !n445 : n445);
assign n792  = /* LUT    2  9  7 */ n76;
assign n793  = /* LUT   11  7  4 */ n541;
assign n794  = /* LUT    4  6  3 */ (n13 ? n20 : 1'b0);
assign n795  = /* LUT    5  5  2 */ (n159 ? (n10 ? 1'b1 : (n11 ? 1'b1 : n49)) : 1'b0);
assign n796  = /* LUT    7  5  4 */ (n4 ? (n22 ? 1'b1 : n63) : 1'b0);
assign n797  = /* LUT    6 12  0 */ (n215 ? (n25 ? (n68 ? !n296 : 1'b1) : 1'b1) : 1'b0);
assign n798  = /* LUT    4 12  1 */ n211;
assign n799  = /* LUT    8 12  2 */ (n68 ? (n25 ? n475 : n464) : n475);
assign n800  = /* LUT    6  4  5 */ (n243 ? (n149 ? 1'b0 : !n229) : (n149 ? !n150 : (n229 ? !n150 : n150)));
assign n801  = /* LUT    8  4  7 */ (n325 ? (n235 ? 1'b1 : n403) : (n235 ? n249 : (n403 ? n249 : !n249)));
assign n802  = /* LUT   12 10  1 */ n555;
assign n803  = /* LUT    7  6  5 */ (n432 ? (n337 ? (n413 ? 1'b1 : !n59) : (n413 ? !n59 : 1'b1)) : (n337 ? (n413 ? 1'b0 : n59) : (n413 ? n59 : 1'b0)));
assign n804  = /* LUT    8 13  3 */ (n275 ? (n31 ? !n483 : 1'b1) : (n31 ? n483 : 1'b0));
assign n805  = /* LUT    7  9  1 */ n355;
assign n806  = /* LUT    9  9  3 */ (n70 ? n498 : n491);
assign n807  = /* LUT    2  5  5 */ (n92 ? !n19 : n19);
assign n808  = /* LUT    6  5  6 */ (n245 ? 1'b0 : !n69);
assign n809  = /* LUT    7 10  2 */ (n362 ? (n25 ? (n68 ? !n365 : 1'b1) : 1'b1) : 1'b0);
assign n810  = /* LUT    5 13  5 */ n219;
assign n811  = /* LUT    2  9  2 */ n34;
assign n812  = /* LUT    7  2  7 */ (n318 ? (n304 ? (n316 ? !n312 : 1'b0) : (n316 ? 1'b0 : !n312)) : (n304 ? (n316 ? 1'b0 : !n312) : (n316 ? !n312 : 1'b0)));
assign n813  = /* LUT    4  9  4 */ n75;
assign n814  = /* LUT    8  8  0 */ (n28 ? (n441 ? !n444 : n444) : (n441 ? n444 : !n444));
assign n815  = /* LUT    6  8  7 */ (n276 ? (n287 ? !n196 : n196) : (n287 ? n196 : !n196));
assign n816  = /* LUT    7 13  3 */ (n25 ? (n68 ? n380 : n43) : n380);
assign n817  = /* LUT    9 13  5 */ n519;
assign n818  = /* LUT    5  5  6 */ (n154 ? (n153 ? 1'b1 : n156) : (n153 ? n157 : (n156 ? n157 : !n157)));
assign n819  = /* LUT    6 12  4 */ (n217 ? (n101 ? (n147 ? !n286 : 1'b1) : (n147 ? 1'b1 : !n286)) : 1'b0);
assign n820  = /* LUT    6  4  0 */ (n246 ? (n232 ? !n237 : n237) : (n232 ? n237 : !n237));
assign n821  = /* LUT    8 12  6 */ n378;
assign n822  = /* LUT    8  4  2 */ (n307 ? (n233 ? n399 : 1'b0) : (n233 ? !n399 : 1'b1));
assign n823  = /* LUT    7  6  0 */ (n37 ? (n334 ? (n327 ? 1'b1 : !n59) : (n327 ? !n59 : 1'b1)) : (n334 ? (n327 ? 1'b0 : n59) : (n327 ? n59 : 1'b0)));
assign n824  = /* LUT    5  9  3 */ n190;
assign n828  = /* LUT    6  5  1 */ (n252 ? (n10 ? 1'b1 : (n11 ? 1'b1 : n49)) : 1'b0);
assign n829  = /* LUT    7  9  5 */ n354;
assign n830  = /* LUT    8  5  3 */ (n253 ? (n170 ? !n18 : 1'b1) : (n170 ? n18 : 1'b0));
assign n831  = /* LUT    9  9  7 */ (n445 ? (n31 ? n500 : 1'b0) : (n31 ? !n500 : 1'b1));
assign n832  = /* LUT    5 12  4 */ n207;
assign n833  = /* LUT    6  8  2 */ (n288 ? (n276 ? (n287 ? !n196 : n196) : (n287 ? n196 : !n196)) : (n276 ? (n287 ? n196 : !n196) : (n287 ? !n196 : n196)));
assign n834  = /* LUT    7 12  6 */ n373;
assign n835  = /* LUT    4  8  3 */ !n73;
assign n836  = /* LUT    8  8  4 */ (n30 ? n436 : !n436);
assign n837  = /* LUT    5  5  1 */ (n250 ? (n10 ? 1'b1 : (n11 ? 1'b1 : n49)) : 1'b0);
assign n838  = /* LUT    7 13  7 */ n384;
assign n839  = /* LUT    7  5  3 */ (n59 ? (n328 ? (n171 ? !n175 : n175) : (n171 ? n175 : !n175)) : 1'b0);
assign n840  = /* LUT    4 12  0 */ n144;
assign n841  = /* LUT    8 12  1 */ (n70 ? !n387 : !n512);
assign n842  = /* LUT    6  4  4 */ (n246 ? (n160 ? !n237 : n237) : (n160 ? n237 : !n237));
assign n843  = /* LUT    8  4  6 */ (n414 ? (n409 ? (n410 ? n416 : !n416) : (n410 ? !n416 : n416)) : (n409 ? (n410 ? !n416 : n416) : (n410 ? n416 : !n416)));
assign n844  = /* LUT   12 10  0 */ n228;
assign n845  = /* LUT    6  7  6 */ (n183 ? 1'b0 : !n184);
assign n846  = /* LUT    7  9  0 */ (n70 ? !n448 : !n450);
assign n847  = /* LUT    9  6  6 */ (n493 ? !n418 : n418);
assign n848  = /* LUT    1  6  6 */ n17;
assign n849  = /* LUT    9  9  2 */ (n445 ? (n442 ? (n501 ? !n31 : 1'b1) : (n501 ? n31 : 1'b0)) : (n442 ? (n501 ? n31 : 1'b0) : (n501 ? !n31 : 1'b1)));
assign n850  = /* LUT   11 11  5 */ n511;
assign n854  = /* LUT    6 11  3 */ n291;
assign n855  = /* LUT    8 11  5 */ n466;
assign n856  = /* LUT    7 12  1 */ n375;
assign n857  = /* LUT    9 12  3 */ (n70 ? n41 : n524);
assign n858  = /* LUT    5  4  4 */ (n106 ? (n10 ? 1'b0 : (n11 ? 1'b0 : !n49)) : 1'b0);
assign n859  = /* LUT    6  8  6 */ (n122 ? (n276 ? n287 : !n287) : (n276 ? !n287 : n287));
assign n860  = /* LUT    7  4  6 */ (n329 ? (n155 ? !n236 : n236) : (n155 ? n236 : !n236));
assign n861  = /* LUT    7 13  2 */ n376;
assign n862  = /* LUT    5  5  5 */ (n180 ? (n10 ? 1'b0 : (n11 ? 1'b0 : !n49)) : 1'b0);
assign n863  = /* LUT    7  5  7 */ (n4 ? (n18 ? !n63 : n22) : 1'b0);
assign n864  = /* LUT    8  4  1 */ (n405 ? (n415 ? (n411 ? !n408 : n408) : (n411 ? n408 : !n408)) : (n415 ? (n411 ? n408 : !n408) : (n411 ? !n408 : n408)));
assign n865  = /* LUT    2  4  7 */ (n10 ? 1'b0 : !n49);
assign n866  = /* LUT    6  7  1 */ (n276 ? (n259 ? n264 : !n264) : (n259 ? !n264 : n264));
assign n867  = /* LUT    8  7  3 */ (n27 ? (n426 ? (n254 ? n434 : !n434) : n434) : (n426 ? n254 : 1'b0));
assign n868  = /* LUT    5  8  6 */ (n182 ? (n163 ? n88 : 1'b1) : (n163 ? !n88 : 1'b0));
assign n869  = /* LUT    9  8  1 */ n497;
assign n870  = /* LUT    5 11  2 */ n198;
assign n871  = /* LUT    4  4  5 */ n106;
assign n872  = /* LUT    7 11  4 */ (n176 ? (n31 ? n465 : 1'b0) : (n31 ? !n465 : 1'b1));
assign n873  = /* LUT    4  7  1 */ n118;
assign n874  = /* LUT    1  3  4 */ (n56 ? (n8 ? 1'b0 : !n51) : (n8 ? !n51 : 1'b0));
assign n875  = /* LUT    8 11  0 */ (n25 ? (n68 ? 1'b1 : !n477) : (n68 ? !n475 : 1'b1));
assign n876  = /* LUT    6 11  7 */ n290;
assign n877  = /* LUT   11  6  7 */ n439;
assign n878  = /* LUT   11  9  3 */ (n70 ? n549 : n554);
assign n879  = /* LUT    5 12  3 */ n209;
assign n880  = /* LUT    7 12  5 */ (n286 ? n464 : (n167 ? n470 : !n470));
assign n881  = /* LUT    6  8  1 */ (n259 ? n264 : !n264);
assign n882  = /* LUT    4  8  2 */ n78;
assign n883  = /* LUT    9 12  7 */ (n275 ? (n31 ? !n87 : 1'b1) : (n31 ? n87 : 1'b0));
assign n884  = /* LUT    8  8  3 */ (n427 ? (n97 ? n274 : !n274) : (n97 ? !n274 : n274));
assign n885  = /* LUT    7  4  1 */ (n307 ? (n415 ? (n326 ? 1'b0 : !n401) : (n326 ? 1'b1 : n401)) : (n415 ? (n326 ? 1'b1 : n401) : (n326 ? 1'b0 : !n401)));
assign n886  = /* LUT    5  5  0 */ (n16 ? (n10 ? 1'b0 : (n11 ? 1'b0 : !n49)) : 1'b0);
assign n887  = /* LUT    7  5  2 */ (n4 ? !n19 : 1'b0);
assign n888  = /* LUT    9  5  4 */ n39;
assign n889  = /* LUT    4 11  3 */ n138;
assign n890  = /* LUT    2  3  6 */ (n56 ? (n8 ? 1'b0 : (n7 ? 1'b0 : !n6)) : 1'b0);
assign n891  = /* LUT    6  7  5 */ (n264 ? (n270 ? !n262 : n262) : (n270 ? n262 : !n262));
assign n892  = /* LUT    8  7  7 */ (n438 ? (n435 ? (n425 ? !n274 : n274) : (n425 ? n274 : !n274)) : (n435 ? (n425 ? n274 : !n274) : (n425 ? !n274 : n274)));
assign n893  = /* LUT    5  8  1 */ n178;
assign n894  = /* LUT    7  8  3 */ (n261 ? (n352 ? (n262 ? !n351 : n351) : n351) : (n352 ? n262 : 1'b1));
assign n895  = /* LUT    4  4  0 */ n113;
assign n896  = /* LUT    9  8  5 */ (n493 ? (n275 ? n418 : !n418) : (n275 ? !n418 : n418));
assign n897  = /* LUT    5 11  6 */ n206;
assign n898  = /* LUT    4  7  5 */ n125;
assign n899  = /* LUT    6 11  2 */ (n25 ? 1'b0 : !n68);
assign n900  = /* LUT    8 11  4 */ (n70 ? n465 : n468);
assign n901  = /* LUT   11  9  7 */ (n70 ? n550 : n548);
assign n902  = /* LUT    7 12  0 */ n374;
assign n903  = /* LUT    5 12  7 */ n294;
assign n904  = /* LUT    9 12  2 */ (n70 ? n523 : n515);
assign n905  = /* LUT    7  4  5 */ (n239 ? (n314 ? n315 : !n315) : (n314 ? !n315 : n315));
assign n906  = /* LUT    8  3  5 */ (n315 ? (n404 ? n161 : 1'b1) : (n404 ? (n161 ? n400 : !n400) : !n400));
assign n907  = /* LUT    5  7  4 */ n163;
assign n908  = /* LUT    2  3  1 */ (n54 ? (n48 ? 1'b0 : (n52 ? 1'b1 : !n9)) : 1'b0);
assign n909  = /* LUT    4 11  7 */ n145;
assign n910  = /* LUT    7  7  6 */ (n266 ? (n254 ? n261 : !n261) : (n254 ? !n261 : n261));
assign n911  = /* LUT    4 14  3 */ n45;
assign n912  = /* LUT    8  7  2 */ (n435 ? (n349 ? (n425 ? !n274 : n274) : (n425 ? n274 : !n274)) : (n349 ? (n425 ? n274 : !n274) : (n425 ? !n274 : n274)));
assign n913  = /* LUT   11  5  5 */ n114;
assign n914  = /* LUT    5  8  5 */ n179;
assign n915  = /* LUT    9  8  0 */ n495;
assign n916  = /* LUT    7  8  7 */ (n193 ? (n339 ? 1'b0 : !n255) : (n339 ? 1'b1 : n346));
assign n917  = /* LUT    5 11  1 */ n202;
assign n918  = /* LUT    4  4  4 */ n105;
assign n919  = /* LUT    7 11  3 */ n370;
assign n920  = /* LUT    4  7  0 */ (n119 ? (n28 ? n110 : !n110) : (n28 ? !n110 : n110));
assign n921  = /* LUT    1  3  3 */ (n58 ? (n7 ? 1'b0 : !n51) : (n7 ? !n51 : 1'b0));
assign n922  = /* LUT    2  7  7 */ n73;
assign n923  = /* LUT   11  9  2 */ (n442 ? !n96 : n96);
assign n924  = /* LUT    5 12  2 */ (n286 ? n221 : (n101 ? n147 : !n147));
assign n925  = /* LUT    4  8  1 */ n131;
assign n926  = /* LUT    9 12  6 */ (n176 ? (n31 ? n387 : 1'b0) : (n31 ? !n387 : 1'b1));
assign n927  = /* LUT    7  4  0 */ (n160 ? (n155 ? !n236 : n236) : (n155 ? n236 : !n236));
assign n928  = /* LUT    2 11  4 */ n99;
assign n929  = /* LUT   12 11  7 */ n558;
assign n930  = /* LUT    8  3  0 */ (n161 ? (n404 ? !n315 : 1'b0) : (n404 ? (n315 ? n402 : !n402) : !n402));
assign n931  = /* LUT    6  3  7 */ n228;
assign n932  = /* LUT    4 11  2 */ n204;
assign n933  = /* LUT    7  7  1 */ (n27 ? (n347 ? (n183 ? n184 : 1'b0) : (n183 ? !n184 : 1'b1)) : (n183 ? n184 : 1'b0));
assign n934  = /* LUT    2  3  5 */ (n56 ? (n8 ? (n7 ? 1'b0 : !n6) : 1'b0) : 1'b0);
assign n935  = /* LUT    6  7  4 */ (n264 ? n270 : !n270);
assign n936  = /* LUT    8  7  6 */ (n347 ? (n426 ? n276 : 1'b1) : (n426 ? (n276 ? n434 : !n434) : !n434));
assign n937  = /* LUT    5  8  0 */ n177;
assign n938  = /* LUT    7  8  2 */ (n192 ? (n352 ? (n260 ? n348 : !n348) : !n348) : (n352 ? n260 : 1'b1));
assign n939  = /* LUT   12 12  7 */ n516;
assign n940  = /* LUT    9  8  4 */ n494;
assign n941  = /* LUT    5 11  5 */ (n68 ? (n25 ? n201 : n194) : n201);
assign n942  = /* LUT    7 11  7 */ (n28 ? (n31 ? !n369 : 1'b1) : (n31 ? n369 : 1'b0));
assign n943  = /* LUT    4  7  4 */ (n121 ? (n119 ? (n110 ? 1'b1 : n88) : (n110 ? n88 : 1'b1)) : (n119 ? (n110 ? 1'b0 : !n88) : (n110 ? !n88 : 1'b0)));
assign n944  = /* LUT   11  6  1 */ n490;
assign n945  = /* LUT    5 14  7 */ n224;
assign n946  = /* LUT    6 10  5 */ n280;
assign n947  = /* LUT   11  9  6 */ (n440 ? (n31 ? !n550 : 1'b1) : (n31 ? n550 : 1'b0));
assign n948  = /* LUT    8 10  7 */ (n28 ? (n445 ? (n459 ? !n31 : 1'b1) : (n459 ? n31 : 1'b0)) : (n445 ? (n459 ? n31 : 1'b0) : (n459 ? !n31 : 1'b1)));
assign n949  = /* LUT    6 13  1 */ n300;
assign n950  = /* LUT    8  2  3 */ (n312 ? (n308 ? (n398 ? 1'b1 : n306) : (n398 ? n306 : 1'b1)) : (n308 ? 1'b0 : n306));
assign n951  = /* LUT    9 11  5 */ n86;
assign n952  = /* LUT   12 11  2 */ n556;
assign n953  = /* LUT    5  6  2 */ (select ? !n164 : 1'b0);
assign n954  = /* LUT    4 10  5 */ n107;
assign n955  = /* LUT    6  3  2 */ (n238 ? (n10 ? 1'b0 : (n11 ? 1'b0 : !n49)) : 1'b0);
assign n956  = /* LUT    8  3  4 */ (n305 ? (n227 ? 1'b1 : n401) : (n227 ? 1'b0 : !n401));
assign n957  = /* LUT   11 12  7 */ (n471 ? (n275 ? (n511 ? !n31 : 1'b1) : (n511 ? n31 : 1'b0)) : (n275 ? (n511 ? n31 : 1'b0) : (n511 ? !n31 : 1'b1)));
assign n958  = /* LUT    2  3  0 */ (n56 ? (n8 ? (n6 ? !n7 : 1'b0) : 1'b0) : 1'b0);
assign n959  = /* LUT    7  7  5 */ (n345 ? (n344 ? n258 : !n258) : (n344 ? !n258 : n258));
assign n960  = /* LUT    4  3  2 */ (n60 ? (n12 ? !rst : 1'b0) : 1'b0);
assign n961  = /* LUT    8  7  1 */ (n193 ? (n255 ? (n346 ? 1'b0 : n339) : n346) : (n255 ? (n346 ? 1'b0 : !n339) : 1'b1));
assign n962  = /* LUT   11  5  4 */ n488;
assign n963  = /* LUT    8  6  5 */ (n339 ? (n346 ? !n255 : (n193 ? !n255 : 1'b1)) : (n346 ? 1'b0 : (n193 ? 1'b1 : !n255)));
assign n964  = /* LUT    5 11  0 */ (n25 ? (n68 ? 1'b1 : !n85) : (n68 ? !n201 : 1'b1));
assign n965  = /* LUT    7 11  2 */ (n463 ? (n25 ? (n68 ? !n464 : 1'b1) : 1'b1) : 1'b0);
assign n966  = /* LUT    2  6  1 */ (rst ? 1'b1 : (n67 ? n64 : 1'b0));
assign n967  = /* LUT    5 14  2 */ n225;
assign n968  = /* LUT    6 10  0 */ n283;
assign n969  = /* LUT    7 14  4 */ n391;
assign n970  = /* LUT   11  9  1 */ (n137 ? (n31 ? !n83 : 1'b1) : (n31 ? n83 : 1'b0));
assign n971  = /* LUT    8 10  2 */ (n28 ? (n31 ? !n460 : 1'b1) : (n31 ? n460 : 1'b0));
assign n972  = /* LUT    9 14  6 */ n525;
assign n973  = /* LUT    6 13  5 */ n303;
assign n974  = /* LUT    8  2  7 */ (n398 ? n311 : (n308 ? 1'b1 : n306));
assign n975  = /* LUT    7  3  3 */ (n161 ? (n315 ? (n160 ? n324 : !n324) : n160) : (n315 ? 1'b0 : n324));
assign n976  = /* LUT    4 10  0 */ n140;
assign n977  = /* LUT    2 10  7 */ n81;
assign n978  = /* LUT    5  6  6 */ n16;
assign n979  = /* LUT    6 14  6 */ !n70;
assign n980  = /* LUT    6  3  6 */ (n239 ? n314 : !n314);
assign n981  = /* LUT    4  2  5 */ (n49 ? (n55 ? 1'b0 : (n9 ? !n52 : 1'b1)) : (n9 ? !n52 : 1'b1));
assign n982  = /* LUT    6  6  2 */ n167;
assign n983  = /* LUT    7 15  4 */ n397;
assign n984  = /* LUT    4 11  1 */ n139;
assign n985  = /* LUT    7  7  0 */ (n254 ? (n276 ? (n347 ? 1'b0 : !n27) : (n347 ? !n27 : 1'b0)) : (n276 ? (n347 ? 1'b0 : n27) : (n347 ? n27 : 1'b0)));
assign n986  = /* LUT    2  3  4 */ (n10 ? (n50 ? (n60 ? n12 : 1'b1) : 1'b0) : (n60 ? n12 : 1'b1));
assign n987  = /* LUT    8  6  0 */ (n256 ? (n183 ? (n430 ? !n428 : n428) : !n430) : (n183 ? 1'b0 : !n428));
assign n988  = /* LUT    6  9  3 */ (n269 ? (n24 ? (n353 ? !n286 : 1'b1) : (n353 ? 1'b1 : !n286)) : 1'b0);
assign n989  = /* LUT    8  9  5 */ (n70 ? n449 : n452);
assign n990  = /* LUT    2  6  5 */ (n63 ? (n22 ? n18 : 1'b0) : 1'b0);
assign n991  = /* LUT    5 14  6 */ (n68 ? (n25 ? n220 : n221) : n220);
assign n992  = /* LUT    9 14  1 */ n527;
assign n993  = /* LUT    4  6  7 */ (n119 ? !n110 : n110);
assign n994  = /* LUT    6 10  4 */ n284;
assign n995  = /* LUT    8 10  6 */ (n445 ? (n31 ? n453 : 1'b0) : (n31 ? !n453 : 1'b1));
assign n996  = /* LUT    6 13  0 */ n299;
assign n997  = /* LUT   11  8  0 */ (select ? 1'b1 : n29);
assign n998  = /* LUT    8  2  2 */ (n306 ? (n308 ? (n398 ? 1'b0 : n312) : n398) : (n308 ? (n398 ? 1'b0 : !n312) : 1'b1));
assign n999  = /* LUT    2 10  2 */ n82;
assign n1000 = /* LUT    7  3  7 */ (n233 ? (n239 ? (n235 ? 1'b0 : !n314) : (n235 ? 1'b1 : n314)) : (n235 ? !n314 : 1'b0));
assign n1001 = /* LUT    4 10  4 */ n134;
assign n1002 = /* LUT    8 14  3 */ n481;
assign n1003 = /* LUT   11 12  6 */ (n275 ? (n31 ? !n41 : 1'b1) : (n31 ? n41 : 1'b0));
assign n1004 = /* LUT    8 13  7 */ (n70 ? n482 : n486);
assign n1005 = /* LUT    7  7  4 */ (n260 ? (n262 ? (n192 ? 1'b0 : !n261) : (n192 ? 1'b1 : n261)) : (n192 ? !n261 : 1'b0));
assign n1006 = /* LUT    5 10  4 */ n132;
assign n1007 = /* LUT    5 13  0 */ (n25 ? (n68 ? 1'b1 : !n298) : (n68 ? !n218 : 1'b1));
assign n1008 = /* LUT    7 10  6 */ n279;
assign n1009 = /* LUT    8  6  4 */ (n193 ? (n346 ? (n255 ? n339 : !n339) : (n255 ? 1'b0 : n339)) : (n346 ? (n255 ? !n339 : 1'b0) : 1'b1));
assign n1010 = /* LUT    7  2  2 */ (n317 ? n406 : !n406);
assign n1011 = /* LUT    8  9  0 */ (n176 ? (n437 ? !n445 : n445) : (n437 ? n445 : !n445));
assign n1012 = /* LUT    1  5  2 */ !n13;
assign n1013 = /* LUT    6  9  7 */ (n286 ? n98 : (n24 ? n353 : !n353));
assign n1014 = /* LUT    2  6  0 */ (n13 ? 1'b0 : (n61 ? 1'b0 : (n62 ? 1'b0 : !n20)));
assign n1015 = /* LUT    5 14  1 */ n223;
assign n1016 = /* LUT    4  6  2 */ (n59 ? (n111 ? !n173 : n173) : 1'b0);
assign n1017 = /* LUT    7 14  3 */ n394;
assign n1018 = /* LUT    8 10  1 */ (n28 ? (n176 ? (n214 ? !n31 : 1'b1) : (n214 ? n31 : 1'b0)) : (n176 ? (n214 ? n31 : 1'b0) : (n214 ? !n31 : 1'b1)));
assign n1019 = /* LUT    9 14  5 */ n526;
assign n1020 = /* LUT    6 13  4 */ n302;
assign n1021 = /* LUT    8  2  6 */ (n398 ? (n306 ? (n312 ? n308 : !n308) : n312) : (n306 ? n308 : (n312 ? n308 : !n308)));
assign n1022 = /* LUT   11  8  4 */ n333;
assign n1023 = /* LUT    7  3  2 */ (n314 ? !n235 : 1'b0);
assign n1024 = /* LUT    2 10  6 */ n74;
assign n1025 = /* LUT    5  6  5 */ n162;
assign n1026 = /* LUT   12 11  5 */ n557;
assign n1027 = /* LUT    2  2  2 */ (rst ? 1'b0 : (n48 ? 1'b1 : (n10 ? n50 : 1'b0)));
assign n1028 = /* LUT    7  6  4 */ (n63 ? (n22 ? (n19 ? 1'b1 : n21) : 1'b1) : (n22 ? 1'b1 : (n19 ? n21 : 1'b1)));
assign n1029 = /* LUT   11 12  1 */ (n273 ? (n31 ? n523 : 1'b0) : (n31 ? !n523 : 1'b1));
assign n1030 = /* LUT    8 13  2 */ (n70 ? n479 : n484);
assign n1031 = /* LUT    5  9  7 */ (n68 ? (n25 ? n187 : n98) : n187);
assign n1032 = /* LUT    2  5  4 */ (n91 ? !n63 : n63);
assign n1033 = /* LUT    6  5  5 */ (n245 ? (n242 ? 1'b0 : !n241) : (n242 ? !n69 : (n241 ? !n69 : n69)));
assign n1034 = /* LUT    8  5  7 */ (n407 ? !n416 : n416);
assign n1035 = /* LUT    7 10  1 */ (n70 ? !n453 : !n456);
assign n1036 = /* LUT    5 13  4 */ n210;
assign n1037 = /* LUT    6  9  2 */ (n25 ? (n68 ? 1'b1 : !n188) : (n68 ? !n187 : 1'b1));
assign n1038 = /* LUT    7  2  6 */ (n313 ? (n227 ? (n152 ? 1'b0 : n321) : (n152 ? n321 : 1'b0)) : (n227 ? (n152 ? 1'b1 : !n321) : (n152 ? !n321 : 1'b1)));
assign n1039 = /* LUT    4  9  3 */ (n25 ? (n68 ? n188 : n98) : n188);
assign n1040 = /* LUT    8  9  4 */ (n442 ? (n31 ? !n447 : 1'b1) : (n31 ? n447 : 1'b0));
assign n1041 = /* LUT   11  7  7 */ (n537 ? (n71 ? n88 : 1'b1) : (n71 ? !n88 : 1'b0));
assign n1042 = /* LUT    4  6  6 */ (select ? !n116 : 1'b0);
assign n1043 = /* LUT    8  2  1 */ (n398 ? (n312 ? (n306 ? 1'b0 : n308) : n306) : (n312 ? (n306 ? 1'b0 : !n308) : 1'b1));
assign n1044 = /* LUT    6 12  3 */ (n292 ? (n25 ? (n68 ? !n43 : 1'b1) : 1'b1) : 1'b0);
assign n1045 = /* LUT    8 12  5 */ n476;
assign n1046 = /* LUT    5  6  0 */ (n172 ? (n108 ? (n175 ? !n59 : 1'b1) : (n175 ? 1'b1 : !n59)) : (n108 ? (n175 ? n59 : 1'b0) : (n175 ? 1'b0 : n59)));
assign n1047 = /* LUT    5  9  2 */ n186;
assign n1048 = /* LUT    6  5  0 */ (n333 ? (n10 ? 1'b0 : (n11 ? 1'b0 : !n49)) : 1'b0);
assign n1049 = /* LUT    8 13  6 */ (n446 ? (n31 ? !n479 : 1'b1) : (n31 ? n479 : 1'b0));
assign n1050 = /* LUT    4  5  1 */ (n13 ? !n20 : n20);
assign n1051 = /* LUT    9  9  6 */ (n70 ? n500 : n499);
assign n1052 = /* LUT    7  9  4 */ n189;
assign n1053 = /* LUT    8  5  2 */ (n253 ? (n408 ? (n332 ? n335 : 1'b1) : (n332 ? !n335 : 1'b0)) : (n408 ? (n332 ? !n335 : 1'b0) : (n332 ? n335 : 1'b1)));
assign n1054 = /* LUT   11  3  5 */ n533;
assign n1055 = /* LUT    5 10  3 */ n197;
assign n1056 = /* LUT    7 10  5 */ (n286 ? n365 : (n228 ? n462 : !n462));
assign n1057 = /* LUT    8  6  3 */ (n256 ? (n183 ? n428 : (n430 ? n428 : !n428)) : (n183 ? 1'b1 : n430));
assign n1058 = /* LUT    7  2  1 */ (n226 ? 1'b0 : (n309 ? 1'b0 : (n306 ? n311 : 1'b1)));
assign n1059 = /* LUT    6  9  6 */ n272;
assign n1060 = /* LUT    4  9  7 */ n127;
assign n1061 = /* LUT   11  7  2 */ n540;
assign n1062 = /* LUT    5 14  0 */ n46;
assign n1063 = /* LUT    4  6  1 */ (n21 ? !n22 : 1'b0);
assign n1064 = /* LUT    7 14  2 */ (n25 ? (n68 ? n392 : n395) : n392);
assign n1065 = /* LUT    9 14  4 */ n520;
assign n1066 = /* LUT    7 13  6 */ n382;
assign n1067 = /* LUT   11  8  3 */ n545;
assign n1068 = /* LUT    8 12  0 */ (n176 ? n273 : !n273);
assign n1069 = /* LUT    6 12  7 */ n289;
assign n1070 = /* LUT    6  4  3 */ (n14 ? (n10 ? 1'b0 : (n11 ? 1'b0 : !n49)) : 1'b0);
assign n1071 = /* LUT    8  4  5 */ (n248 ? (n314 ? n249 : 1'b1) : (n403 ? (n314 ? 1'b1 : n249) : (n314 ? 1'b0 : !n249)));
assign n1072 = /* LUT    7  6  3 */ (n63 ? !n19 : 1'b0);
assign n1073 = /* LUT    8 13  1 */ (n446 ? (n31 ? !n482 : 1'b1) : (n31 ? n482 : 1'b0));
assign n1074 = /* LUT    5  9  6 */ n185;
assign n1075 = /* LUT    9  9  1 */ (n70 ? !n503 : !n502);
assign n1076 = /* LUT    2  5  3 */ (n90 ? !n62 : n62);
assign n1077 = /* LUT    6  5  4 */ (n251 ? (n10 ? 1'b1 : (n11 ? 1'b1 : n49)) : 1'b0);
assign n1078 = /* LUT   11 11  4 */ n214;
assign n1079 = /* LUT    8  5  6 */ (n411 ? n424 : !n424);
assign n1080 = /* LUT    7 10  0 */ (n389 ? (n340 ? (n372 ? !n286 : 1'b1) : (n372 ? 1'b1 : !n286)) : 1'b0);
assign n1081 = /* LUT    5 10  7 */ (n286 ? n194 : (n148 ? n38 : !n38));
assign n1082 = /* LUT    5 13  3 */ n212;
assign n1083 = /* LUT    2  9  0 */ n36;
assign n1084 = /* LUT    7  2  5 */ (n317 ? (n310 ? (n406 ? 1'b0 : !n312) : 1'b0) : (n310 ? 1'b0 : (n406 ? !n312 : 1'b0)));
assign n1085 = /* LUT    4  9  2 */ n40;
assign n1086 = /* LUT    8  9  3 */ (n442 ? (n31 ? !n449 : 1'b1) : (n31 ? n449 : 1'b0));
assign n1087 = /* LUT    6  8  5 */ (n268 ? (n276 ? (n287 ? !n196 : n196) : (n287 ? n196 : !n196)) : (n276 ? (n287 ? n196 : !n196) : (n287 ? !n196 : n196)));
assign n1088 = /* LUT    8  8  7 */ (n30 ? (n436 ? (n97 ? n274 : !n274) : (n97 ? !n274 : n274)) : (n436 ? (n97 ? !n274 : n274) : (n97 ? n274 : !n274)));
assign n1089 = /* LUT    9 13  3 */ n521;
assign n1090 = /* LUT    5  5  4 */ (n165 ? (n10 ? 1'b0 : (n11 ? 1'b0 : !n49)) : 1'b0);
assign n1091 = /* LUT    6 12  2 */ (n25 ? (n68 ? 1'b1 : !n380) : (n68 ? !n295 : 1'b1));
assign n1092 = /* LUT    7  5  6 */ (n175 ? (n323 ? !n413 : n413) : (n323 ? n413 : !n413));
assign n1093 = /* LUT    8 12  4 */ n473;
assign n1094 = /* LUT    8  4  0 */ (n409 ? !n410 : n410);
assign n1095 = /* LUT    6  4  7 */ (n243 ? 1'b0 : !n150);
assign n1096 = /* LUT    7  6  7 */ n24;
assign n1097 = /* LUT    5  9  1 */ n271;
assign n1098 = /* LUT    7  9  3 */ n357;
assign n1099 = /* LUT    4  5  0 */ (n19 ? 1'b0 : !n21);
assign n1100 = /* LUT    9  9  5 */ (n442 ? (n31 ? !n503 : 1'b1) : (n31 ? n503 : 1'b0));
assign n1101 = /* LUT    2  5  7 */ (n94 ? !n22 : n22);
assign n1102 = /* LUT    8  5  1 */ (n95 ? (n422 ? (n424 ? 1'b1 : !n59) : (n424 ? !n59 : 1'b1)) : (n422 ? (n424 ? 1'b0 : n59) : (n424 ? n59 : 1'b0)));
assign n1103 = /* LUT    7  2  0 */ (n321 ? (n227 ? !n152 : n152) : 1'b0);
assign n1104 = /* LUT   11  7  1 */ (n445 ? n71 : !n71);
assign n1105 = /* LUT    8  8  2 */ (n28 ? !n441 : n441);
assign n1106 = /* LUT    7 13  5 */ n381;
assign n1107 = /* LUT    7  5  1 */ (n244 ? !n417 : !n338);
assign n1108 = /* LUT    9 13  7 */ n340;
assign n1109 = /* LUT    6 12  6 */ (n68 ? (n25 ? n295 : n43) : n295);
assign n1110 = /* LUT    6  4  2 */ (n247 ? (n232 ? (n158 ? !n237 : n237) : (n158 ? n237 : !n237)) : (n232 ? (n158 ? n237 : !n237) : (n158 ? !n237 : n237)));
assign n1111 = /* LUT    8  4  4 */ (n248 ? (n314 ? n403 : 1'b1) : (n314 ? (n403 ? n249 : !n249) : n249));
assign n1112 = /* LUT    7  6  2 */ (n4 ? !n336 : 1'b0);
assign n1113 = /* LUT    9  9  0 */ (n70 ? !n83 : !n506);
assign n1114 = /* LUT    2  5  2 */ (n89 ? !n61 : n61);
assign n1115 = /* LUT   11 11  3 */ (n100 ? !n421 : n421);
assign n1116 = /* LUT    6 11  1 */ (n285 ? (n168 ? (n366 ? !n286 : 1'b1) : (n366 ? 1'b1 : !n286)) : 1'b0);
assign n1117 = /* LUT    8 11  3 */ n469;
assign n58   = /* CARRY  1  3  2 */ (1'b0 & n6) | ((1'b0 | n6) & n57);
assign n57   = /* CARRY  1  3  1 */ (1'b0 & n8) | ((1'b0 | n8) & n560);
assign n94   = /* CARRY  2  5  6 */ (1'b0 & n21) | ((1'b0 | n21) & n93);
assign n89   = /* CARRY  2  5  1 */ (1'b0 & n20) | ((1'b0 | n20) & n559);
assign n93   = /* CARRY  2  5  5 */ (1'b0 & n19) | ((1'b0 | n19) & n92);
assign n559  = /* CARRY  2  5  0 */ (n13 & 1'b0) | ((n13 | 1'b0) & n827);
assign n560  = /* CARRY  1  3  0 */ (n56 & 1'b0) | ((n56 | 1'b0) & n853);
assign n92   = /* CARRY  2  5  4 */ (1'b0 & n63) | ((1'b0 | n63) & n91);
assign n91   = /* CARRY  2  5  3 */ (1'b0 & n62) | ((1'b0 | n62) & n90);
assign n90   = /* CARRY  2  5  2 */ (1'b0 & n61) | ((1'b0 | n61) & n89);
/* FF  5 12  6 */ always @(posedge clk) if (1'b1) n212 <= 1'b0 ? 1'b0 : n561;
/* FF  9 12  1 */ always @(posedge clk) if (1'b1) n511 <= 1'b0 ? 1'b0 : n562;
/* FF  2  8  3 */ always @(posedge clk) if (n65) d_vld <= 1'b0 ? 1'b0 : n563;
/* FF  6  8  4 */ assign n263 = n564;
/* FF  4  8  5 */ always @(posedge clk) if (1'b1) n126 <= 1'b0 ? 1'b0 : n565;
/* FF  8  8  6 */ assign n275 = n566;
/* FF  7  4  4 */ assign n324 = n567;
/* FF  1  7  4 */ always @(posedge clk) if (1'b1) n23 <= n1 ? 1'b1 : n568;
/* FF  7 13  0 */ always @(posedge clk) if (1'b1) n381 <= 1'b0 ? 1'b0 : n569;
/* FF  9 13  2 */ always @(posedge clk) if (1'b1) n519 <= 1'b0 ? 1'b0 : n570;
/* FF  5  5  3 */ assign n155 = n571;
/* FF  7  5  5 */ assign n332 = n572;
/* FF  4 12  2 */ always @(posedge clk) if (1'b1) n144 <= 1'b0 ? 1'b0 : n573;
/* FF  8 12  3 */ always @(posedge clk) if (1'b1) n473 <= 1'b0 ? 1'b0 : n574;
/* FF  9  5  7 */ always @(posedge clk) if (1'b1) n489 <= 1'b0 ? 1'b0 : n575;
/* FF  6  4  6 */ assign n160 = n576;
/* FF  5  9  0 */ always @(posedge clk) if (1'b1) n185 <= 1'b0 ? 1'b0 : n577;
/* FF  7  9  2 */ always @(posedge clk) if (1'b1) n355 <= 1'b0 ? 1'b0 : n578;
/* FF  9  9  4 */ always @(posedge clk) if (1'b1) n500 <= 1'b0 ? 1'b0 : n579;
/* FF  5  8  4 */ always @(posedge clk) if (1'b1) n179 <= 1'b0 ? 1'b0 : n580;
/* FF  7  8  6 */ assign n351 = n581;
/* FF  1  3  2 */ always @(posedge clk) if (n53) n6 <= rst ? 1'b0 : n582;
/* FF  8 11  7 */ always @(posedge clk) if (1'b1) n469 <= 1'b0 ? 1'b0 : n583;
/* FF 11  6  5 */ always @(posedge clk) if (1'b1) n417 <= 1'b0 ? 1'b0 : n584;
/* FF  5 12  1 */ always @(posedge clk) if (1'b1) n208 <= 1'b0 ? 1'b0 : n585;
/* FF  7 12  3 */ always @(posedge clk) if (1'b1) n376 <= 1'b0 ? 1'b0 : n586;
/* FF  9 12  5 */ always @(posedge clk) if (1'b1) n515 <= 1'b0 ? 1'b0 : n587;
/* FF  8  8  1 */ assign n441 = n588;
/* FF  7 13  4 */ always @(posedge clk) if (1'b1) n384 <= 1'b0 ? 1'b0 : n589;
/* FF  7  5  0 */ assign n328 = n590;
/* FF  9 13  6 */ always @(posedge clk) if (1'b1) n521 <= 1'b0 ? 1'b0 : n591;
/* FF  5  5  7 */ always @(posedge clk) if (n4) n159 <= 1'b0 ? 1'b0 : n592;
/* FF  9  5  2 */ always @(posedge clk) if (1'b1) n114 <= 1'b0 ? 1'b0 : n593;
/* FF 12  9  5 */ always @(posedge clk) if (1'b1) n554 <= n3 ? 1'b1 : n594;
/* FF  4 12  6 */ always @(posedge clk) if (1'b1) n145 <= 1'b0 ? 1'b0 : n595;
/* FF  8  4  3 */ assign n173 = n596;
/* FF  6  7  3 */ assign n256 = n597;
/* FF  8  7  5 */ assign n437 = n598;
/* FF  7  8  1 */ assign n97 = n599;
/* FF  9  8  3 */ always @(posedge clk) if (1'b1) n495 <= 1'b0 ? 1'b0 : n600;
/* FF  5 11  4 */ always @(posedge clk) if (1'b1) n194 <= 1'b0 ? 1'b0 : n601;
/* FF  7 11  6 */ always @(posedge clk) if (1'b1) n371 <= 1'b0 ? 1'b0 : n602;
/* FF  4  7  3 */ always @(posedge clk) if (1'b1) n119 <= 1'b0 ? 1'b0 : n603;
/* FF  6 11  0 */ assign n287 = n604;
/* FF 11  6  0 */ assign \d_out[5]  = n605;
/* FF  8 11  2 */ always @(posedge clk) if (1'b1) n465 <= 1'b0 ? 1'b0 : n606;
/* FF 11  9  5 */ always @(posedge clk) if (1'b1) n550 <= 1'b0 ? 1'b0 : n607;
/* FF  9 12  0 */ assign n462 = n608;
/* FF  6  8  3 */ assign n262 = n609;
/* FF  7 12  7 */ always @(posedge clk) if (1'b1) n378 <= 1'b0 ? 1'b0 : n610;
/* FF  4  8  4 */ always @(posedge clk) if (1'b1) n125 <= 1'b0 ? 1'b0 : n611;
/* FF  7  4  3 */ assign n314 = n612;
/* FF  8  8  5 */ assign n445 = n613;
/* FF 11 10  6 */ always @(posedge clk) if (1'b1) n552 <= n1 ? 1'b1 : n614;
/* FF  8  3  3 */ assign n407 = n615;
/* FF  6  6  6 */ always @(posedge clk) if (n4) n252 <= 1'b0 ? 1'b0 : n616;
/* FF  8  7  0 */ assign n433 = n617;
/* FF  6  7  7 */ assign n184 = n618;
/* FF 11 13  7 */ always @(posedge clk) if (1'b1) n530 <= 1'b0 ? 1'b0 : n619;
/* FF 11  5  3 */ always @(posedge clk) if (1'b1) n14 <= 1'b0 ? 1'b0 : n620;
/* FF  1  6  7 */ always @(posedge clk) if (1'b1) n17 <= 1'b0 ? 1'b0 : n621;
/* FF  5  8  3 */ always @(posedge clk) if (1'b1) n148 <= 1'b0 ? 1'b0 : n622;
/* FF  7  8  5 */ assign n341 = n623;
/* FF  7 11  1 */ assign n359 = n624;
/* FF  9  8  7 */ always @(posedge clk) if (1'b1) n497 <= 1'b0 ? 1'b0 : n625;
/* FF  1  3  1 */ assign n626 = n627;
/* FF  6 11  4 */ always @(posedge clk) if (1'b1) n290 <= 1'b0 ? 1'b0 : n628;
/* FF 11  6  4 */ always @(posedge clk) if (1'b1) n24 <= 1'b0 ? 1'b0 : n629;
/* FF  8 11  6 */ always @(posedge clk) if (1'b1) n468 <= 1'b0 ? 1'b0 : n630;
/* FF 11  9  0 */ assign \d_out[4]  = n631;
/* FF  5 12  0 */ always @(posedge clk) if (1'b1) n207 <= 1'b0 ? 1'b0 : n632;
/* FF  7 12  2 */ always @(posedge clk) if (1'b1) n375 <= 1'b0 ? 1'b0 : n633;
/* FF  9 12  4 */ always @(posedge clk) if (1'b1) n514 <= 1'b0 ? 1'b0 : n634;
/* FF  5  4  5 */ always @(posedge clk) if (n4) n151 <= 1'b0 ? 1'b0 : n635;
/* FF  7  4  7 */ assign n248 = n636;
/* FF 11 10  1 */ assign \d_out[2]  = n637;
/* FF  6  6  1 */ always @(posedge clk) if (n4) n240 <= 1'b0 ? 1'b0 : n638;
/* FF  8  3  7 */ assign n410 = n639;
/* FF  4 11  0 */ always @(posedge clk) if (1'b1) n138 <= 1'b0 ? 1'b0 : n640;
/* FF  2  3  3 */ assign n53 = n641;
/* FF  2 14  3 */ always @(posedge clk) if (1'b1) n45 <= 1'b0 ? 1'b0 : n642;
/* FF  4  3  5 */ always @(posedge clk) if (1'b1) n60 <= 1'b0 ? 1'b0 : n643;
/* FF  6  7  2 */ assign n255 = n644;
/* FF  8  7  4 */ assign n436 = n645;
/* FF  7  8  0 */ assign n348 = n646;
/* FF  5  8  7 */ always @(posedge clk) if (1'b1) n182 <= 1'b0 ? 1'b0 : n647;
/* FF  9  8  2 */ always @(posedge clk) if (1'b1) n494 <= 1'b0 ? 1'b0 : n648;
/* FF  5 11  3 */ always @(posedge clk) if (1'b1) n203 <= 1'b0 ? 1'b0 : n649;
/* FF  7 11  5 */ always @(posedge clk) if (1'b1) n370 <= 1'b0 ? 1'b0 : n650;
/* FF  4  7  2 */ always @(posedge clk) if (1'b1) n118 <= 1'b0 ? 1'b0 : n651;
/* FF  8 11  1 */ always @(posedge clk) if (1'b1) n464 <= 1'b0 ? 1'b0 : n652;
/* FF  6 10  3 */ always @(posedge clk) if (1'b1) n280 <= 1'b0 ? 1'b0 : n653;
/* FF 11  9  4 */ always @(posedge clk) if (1'b1) n549 <= 1'b0 ? 1'b0 : n654;
/* FF  8 10  5 */ always @(posedge clk) if (1'b1) n458 <= 1'b0 ? 1'b0 : n655;
/* FF  5  4  0 */ assign n149 = n656;
/* FF  7  4  2 */ assign n315 = n657;
/* FF  9 11  3 */ always @(posedge clk) if (1'b1) n100 <= 1'b0 ? 1'b0 : n658;
/* FF  2 10  1 */ always @(posedge clk) if (1'b1) n78 <= 1'b0 ? 1'b0 : n659;
/* FF  7  3  6 */ assign n312 = n660;
/* FF  6  3  0 */ assign n227 = n661;
/* FF  8  3  2 */ assign n405 = n662;
/* FF  2  2  6 */ always @(posedge clk) if (1'b1) n9 <= 1'b0 ? 1'b0 : n663;
/* FF  6  6  5 */ always @(posedge clk) if (n4) n250 <= 1'b0 ? 1'b0 : n664;
/* FF  9  4  0 */ always @(posedge clk) if (1'b1) n228 <= 1'b0 ? 1'b0 : n665;
/* FF  7 15  7 */ always @(posedge clk) if (1'b1) n397 <= 1'b0 ? 1'b0 : n666;
/* FF  4 11  4 */ always @(posedge clk) if (1'b1) n77 <= 1'b0 ? 1'b0 : n667;
/* FF  7  7  3 */ assign n344 = n668;
/* FF  4  3  0 */ assign n88 = n669;
/* FF  9  7  5 */ always @(posedge clk) if (1'b1) n491 <= n3 ? 1'b0 : n670;
/* FF  2  3  7 */ always @(posedge clk) if (n53) n56 <= rst ? 1'b0 : n671;
/* FF  5  8  2 */ always @(posedge clk) if (1'b1) n178 <= 1'b0 ? 1'b0 : n672;
/* FF  7  8  4 */ assign n30 = n673;
/* FF  7 11  0 */ assign n366 = n674;
/* FF  5 11  7 */ always @(posedge clk) if (1'b1) n206 <= 1'b0 ? 1'b0 : n675;
/* FF  8 10  0 */ always @(posedge clk) if (1'b1) n453 <= 1'b0 ? 1'b0 : n676;
/* FF  6 10  7 */ always @(posedge clk) if (1'b1) n284 <= 1'b0 ? 1'b0 : n677;
/* FF  6 13  3 */ always @(posedge clk) if (1'b1) n299 <= 1'b0 ? 1'b0 : n678;
/* FF  8  2  5 */ assign n249 = n679;
/* FF  9 11  7 */ always @(posedge clk) if (1'b1) n510 <= 1'b0 ? 1'b0 : n680;
/* FF  7  3  1 */ assign n317 = n681;
/* FF  9  3  3 */ always @(posedge clk) if (1'b1) n238 <= 1'b0 ? 1'b0 : n682;
/* FF  5  6  4 */ always @(posedge clk) if (1'b1) n165 <= 1'b0 ? 1'b0 : n683;
/* FF  2  2  1 */ assign n48 = n684;
/* FF  6  3  4 */ assign n230 = n685;
/* FF  4 10  7 */ always @(posedge clk) if (1'b1) n136 <= 1'b0 ? 1'b0 : n686;
/* FF  8  3  6 */ assign n171 = n687;
/* FF 11 12  0 */ always @(posedge clk) if (1'b1) n485 <= 1'b0 ? 1'b0 : n688;
/* FF  7 15  2 */ always @(posedge clk) if (1'b1) n395 <= 1'b0 ? 1'b0 : n689;
/* FF 11  4  5 */ always @(posedge clk) if (1'b1) n533 <= n1 ? 1'b1 : n690;
/* FF  5  7  5 */ always @(posedge clk) if (1'b1) n174 <= n1 ? 1'b0 : n691;
/* FF  2  3  2 */ assign n52 = n692;
/* FF  7  7  7 */ assign n193 = n693;
/* FF  8  6  7 */ assign n431 = n694;
/* FF  6  9  1 */ assign n259 = n695;
/* FF  2  6  3 */ assign n66 = n696;
/* FF  5 14  4 */ always @(posedge clk) if (1'b1) n47 <= 1'b0 ? 1'b0 : n697;
/* FF  6 10  2 */ always @(posedge clk) if (1'b1) n279 <= 1'b0 ? 1'b0 : n698;
/* FF  7 14  6 */ always @(posedge clk) if (1'b1) n394 <= 1'b0 ? 1'b0 : n699;
/* FF  8 10  4 */ always @(posedge clk) if (1'b1) n457 <= 1'b0 ? 1'b0 : n700;
/* FF  8  2  0 */ assign n398 = n701;
/* FF  6 13  7 */ always @(posedge clk) if (1'b1) n303 <= 1'b0 ? 1'b0 : n702;
/* FF  6  2  7 */ assign n226 = n703;
/* FF 11  8  7 */ always @(posedge clk) if (1'b1) n545 <= 1'b0 ? 1'b0 : n704;
/* FF  9 11  2 */ always @(posedge clk) if (1'b1) n508 <= 1'b0 ? 1'b0 : n705;
/* FF  2 10  0 */ always @(posedge clk) if (1'b1) n40 <= 1'b0 ? 1'b0 : n706;
/* FF  7  3  5 */ assign n321 = n707;
/* FF  4 10  2 */ always @(posedge clk) if (1'b1) n132 <= 1'b0 ? 1'b0 : n708;
/* FF  9  3  7 */ always @(posedge clk) if (1'b1) n101 <= 1'b0 ? 1'b0 : n709;
/* FF  8  3  1 */ assign n406 = n710;
/* FF  4  2  7 */ always @(posedge clk) if (1'b1) n4 <= 1'b0 ? 1'b0 : n711;
/* FF  7  7  2 */ assign n339 = n712;
/* FF  5 10  2 */ assign n196 = n713;
/* FF  7 10  4 */ assign n122 = n714;
/* FF 11  5  1 */ always @(posedge clk) if (1'b1) n531 <= 1'b0 ? 1'b0 : n715;
/* FF  8  6  2 */ assign n426 = n716;
/* FF  6  9  5 */ assign n270 = n717;
/* FF  4  9  6 */ always @(posedge clk) if (1'b1) n98 <= 1'b0 ? 1'b0 : n718;
/* FF  8  9  7 */ always @(posedge clk) if (1'b1) n452 <= 1'b0 ? 1'b0 : n719;
/* FF  4  6  0 */ assign n108 = n720;
/* FF  7 14  1 */ assign n389 = n721;
/* FF  2  6  7 */ always @(posedge clk) if (1'b1) n68 <= n9 ? 1'b1 : n722;
/* FF  9 14  3 */ always @(posedge clk) if (1'b1) n526 <= 1'b0 ? 1'b0 : n723;
/* FF  6 10  6 */ always @(posedge clk) if (1'b1) n283 <= 1'b0 ? 1'b0 : n724;
/* FF  6  2  2 */ assign n1 = n725;
/* FF  6 13  2 */ always @(posedge clk) if (1'b1) n298 <= 1'b0 ? 1'b0 : n726;
/* FF 11  8  2 */ always @(posedge clk) if (1'b1) n544 <= 1'b0 ? 1'b0 : n727;
/* FF  8  2  4 */ assign n402 = n728;
/* FF  7  3  0 */ assign n316 = n729;
/* FF  9 11  6 */ always @(posedge clk) if (1'b1) n478 <= 1'b0 ? 1'b0 : n730;
/* FF  2 10  4 */ always @(posedge clk) if (1'b1) n80 <= 1'b0 ? 1'b0 : n731;
/* FF  5  6  3 */ always @(posedge clk) if (1'b1) n164 <= 1'b0 ? 1'b0 : n732;
/* FF  4 10  6 */ always @(posedge clk) if (1'b1) n135 <= 1'b0 ? 1'b0 : n733;
/* FF  8 13  0 */ assign n470 = n734;
/* FF  6  5  3 */ assign n244 = n735;
/* FF  8  5  5 */ assign n422 = n736;
/* FF  5 10  6 */ always @(posedge clk) if (1'b1) n198 <= 1'b0 ? 1'b0 : n737;
/* FF  9 10  1 */ always @(posedge clk) if (1'b1) n504 <= n3 ? 1'b1 : n738;
/* FF  5 13  2 */ assign n217 = n739;
/* FF  6  9  0 */ assign n266 = n740;
/* FF  8  6  6 */ assign n430 = n741;
/* FF  4  9  1 */ always @(posedge clk) if (1'b1) n34 <= 1'b0 ? 1'b0 : n742;
/* FF  8  9  2 */ always @(posedge clk) if (1'b1) n447 <= 1'b0 ? 1'b0 : n743;
/* FF  7  2  4 */ assign n308 = n744;
/* FF 11  7  5 */ always @(posedge clk) if (1'b1) n432 <= 1'b0 ? 1'b0 : n745;
/* FF  2  6  2 */ assign n5 = n746;
/* FF  4  6  4 */ assign n111 = n747;
/* FF  7 14  5 */ always @(posedge clk) if (1'b1) n393 <= 1'b0 ? 1'b0 : n748;
/* FF  6 10  1 */ always @(posedge clk) if (1'b1) n278 <= 1'b0 ? 1'b0 : n749;
/* FF  8 10  3 */ always @(posedge clk) if (1'b1) n456 <= 1'b0 ? 1'b0 : n750;
/* FF  6 13  6 */ always @(posedge clk) if (1'b1) n302 <= 1'b0 ? 1'b0 : n751;
/* FF  9 11  1 */ always @(posedge clk) if (1'b1) n507 <= 1'b0 ? 1'b0 : n752;
/* FF  7  3  4 */ assign n320 = n753;
/* FF  4 10  1 */ always @(posedge clk) if (1'b1) n131 <= 1'b0 ? 1'b0 : n754;
/* FF  5  6  7 */ always @(posedge clk) if (1'b1) n168 <= 1'b0 ? 1'b0 : n755;
/* FF  2  2  4 */ always @(posedge clk) if (1'b1) n10 <= 1'b0 ? 1'b0 : n756;
/* FF  7  6  6 */ assign n337 = n757;
/* FF 11 12  3 */ always @(posedge clk) if (1'b1) n523 <= 1'b0 ? 1'b0 : n758;
/* FF  8 13  4 */ always @(posedge clk) if (1'b1) n482 <= 1'b0 ? 1'b0 : n759;
/* FF  8  5  0 */ assign n418 = n760;
/* FF  2  5  6 */ always @(posedge clk) if (1'b1) n21 <= n5 ? 1'b0 : n761;
/* FF  6  5  7 */ assign n239 = n762;
/* FF  5 10  1 */ assign n195 = n763;
/* FF  7 10  3 */ assign n362 = n764;
/* FF  8  6  1 */ assign n274 = n765;
/* FF  2  9  3 */ always @(posedge clk) if (1'b1) n33 <= 1'b0 ? 1'b0 : n766;
/* FF  6  9  4 */ assign n269 = n767;
/* FF  4  9  5 */ always @(posedge clk) if (1'b1) n129 <= 1'b0 ? 1'b0 : n768;
/* FF  8  9  6 */ always @(posedge clk) if (1'b1) n451 <= 1'b0 ? 1'b0 : n769;
/* FF 11  7  0 */ always @(posedge clk) if (1'b1) n537 <= 1'b0 ? 1'b0 : n770;
/* FF  7 14  0 */ assign n388 = n771;
/* FF  2  6  6 */ always @(posedge clk) if (1'b1) n25 <= n9 ? 1'b1 : n772;
/* FF 11  8  1 */ assign \d_out[0]  = n773;
/* FF  6 12  5 */ always @(posedge clk) if (1'b1) n294 <= 1'b0 ? 1'b0 : n774;
/* FF  6  4  1 */ assign n232 = n775;
/* FF  8 12  7 */ always @(posedge clk) if (1'b1) n477 <= 1'b0 ? 1'b0 : n776;
/* FF  7  6  1 */ assign n96 = n777;
/* FF  9  6  3 */ always @(posedge clk) if (1'b1) n490 <= n1 ? 1'b1 : n778;
/* FF  5  9  4 */ always @(posedge clk) if (1'b1) n189 <= 1'b0 ? 1'b0 : n779;
/* FF  2  5  1 */ assign n780 = n781;
/* FF  6  5  2 */ assign n243 = n782;
/* FF  7  9  6 */ always @(posedge clk) if (1'b1) n358 <= 1'b0 ? 1'b0 : n783;
/* FF 11 11  2 */ assign \d_out[3]  = n784;
/* FF  8  5  4 */ assign n421 = n785;
/* FF  9 10  0 */ always @(posedge clk) if (1'b1) n505 <= n3 ? 1'b0 : n786;
/* FF  5 13  1 */ assign n216 = n787;
/* FF  7 10  7 */ always @(posedge clk) if (1'b1) n364 <= 1'b0 ? 1'b0 : n788;
/* FF  7  2  3 */ assign n307 = n789;
/* FF  4  9  0 */ always @(posedge clk) if (1'b1) n127 <= 1'b0 ? 1'b0 : n790;
/* FF  8  9  1 */ assign n137 = n791;
/* FF  2  9  7 */ always @(posedge clk) if (1'b1) n74 <= 1'b0 ? 1'b0 : n792;
/* FF 11  7  4 */ always @(posedge clk) if (1'b1) n540 <= 1'b0 ? 1'b0 : n793;
/* FF  4  6  3 */ assign n73 = n794;
/* FF  5  5  2 */ assign n154 = n795;
/* FF  7  5  4 */ assign n170 = n796;
/* FF  6 12  0 */ assign n285 = n797;
/* FF  4 12  1 */ always @(posedge clk) if (1'b1) n143 <= 1'b0 ? 1'b0 : n798;
/* FF  8 12  2 */ always @(posedge clk) if (1'b1) n472 <= 1'b0 ? 1'b0 : n799;
/* FF  6  4  5 */ assign n236 = n800;
/* FF  8  4  7 */ assign n411 = n801;
/* FF 12 10  1 */ always @(posedge clk) if (1'b1) n556 <= 1'b0 ? 1'b0 : n802;
/* FF  7  6  5 */ assign n71 = n803;
/* FF  8 13  3 */ always @(posedge clk) if (1'b1) n481 <= 1'b0 ? 1'b0 : n804;
/* FF  7  9  1 */ always @(posedge clk) if (1'b1) n354 <= 1'b0 ? 1'b0 : n805;
/* FF  9  9  3 */ always @(posedge clk) if (1'b1) n499 <= 1'b0 ? 1'b0 : n806;
/* FF  2  5  5 */ always @(posedge clk) if (1'b1) n19 <= n5 ? 1'b0 : n807;
/* FF  6  5  6 */ assign n247 = n808;
/* FF  7 10  2 */ assign n361 = n809;
/* FF  5 13  5 */ always @(posedge clk) if (1'b1) n220 <= 1'b0 ? 1'b0 : n810;
/* FF  2  9  2 */ always @(posedge clk) if (1'b1) n76 <= 1'b0 ? 1'b0 : n811;
/* FF  7  2  7 */ assign n311 = n812;
/* FF  4  9  4 */ always @(posedge clk) if (1'b1) n128 <= 1'b0 ? 1'b0 : n813;
/* FF  8  8  0 */ assign n440 = n814;
/* FF  6  8  7 */ assign n192 = n815;
/* FF  7 13  3 */ always @(posedge clk) if (1'b1) n383 <= 1'b0 ? 1'b0 : n816;
/* FF  9 13  5 */ always @(posedge clk) if (1'b1) n43 <= 1'b0 ? 1'b0 : n817;
/* FF  5  5  6 */ assign n158 = n818;
/* FF  6 12  4 */ assign n276 = n819;
/* FF  6  4  0 */ assign n161 = n820;
/* FF  8 12  6 */ always @(posedge clk) if (1'b1) n476 <= 1'b0 ? 1'b0 : n821;
/* FF  8  4  2 */ assign n414 = n822;
/* FF  7  6  0 */ assign n72 = n823;
/* FF  5  9  3 */ always @(posedge clk) if (1'b1) n188 <= 1'b0 ? 1'b0 : n824;
/* FF  2  5  0 */ assign n825 = n826;
/* FF  6  5  1 */ assign n242 = n828;
/* FF  7  9  5 */ always @(posedge clk) if (1'b1) n357 <= 1'b0 ? 1'b0 : n829;
/* FF  8  5  3 */ assign n420 = n830;
/* FF  9  9  7 */ always @(posedge clk) if (1'b1) n503 <= 1'b0 ? 1'b0 : n831;
/* FF  5 12  4 */ always @(posedge clk) if (1'b1) n211 <= 1'b0 ? 1'b0 : n832;
/* FF  6  8  2 */ assign n261 = n833;
/* FF  7 12  6 */ always @(posedge clk) if (1'b1) n365 <= 1'b0 ? 1'b0 : n834;
/* FF  4  8  3 */ always @(posedge clk) if (1'b1) n31 <= 1'b0 ? 1'b0 : n835;
/* FF  8  8  4 */ assign n444 = n836;
/* FF  5  5  1 */ assign n153 = n837;
/* FF  7 13  7 */ always @(posedge clk) if (1'b1) n386 <= 1'b0 ? 1'b0 : n838;
/* FF  7  5  3 */ assign n331 = n839;
/* FF  4 12  0 */ always @(posedge clk) if (1'b1) n142 <= 1'b0 ? 1'b0 : n840;
/* FF  8 12  1 */ assign n147 = n841;
/* FF  6  4  4 */ assign n235 = n842;
/* FF  8  4  6 */ assign n175 = n843;
/* FF 12 10  0 */ always @(posedge clk) if (1'b1) n555 <= 1'b0 ? 1'b0 : n844;
/* FF  6  7  6 */ assign n258 = n845;
/* FF  7  9  0 */ assign n353 = n846;
/* FF  9  6  6 */ always @(posedge clk) if (1'b1) n439 <= n1 ? 1'b1 : n847;
/* FF  1  6  6 */ always @(posedge clk) if (1'b1) n16 <= 1'b0 ? 1'b0 : n848;
/* FF  9  9  2 */ always @(posedge clk) if (1'b1) n498 <= 1'b0 ? 1'b0 : n849;
/* FF 11 11  5 */ always @(posedge clk) if (1'b1) n524 <= n3 ? 1'b1 : n850;
/* FF  1  3  0 */ assign n851 = n852;
/* FF  6 11  3 */ always @(posedge clk) if (1'b1) n289 <= 1'b0 ? 1'b0 : n854;
/* FF  8 11  5 */ always @(posedge clk) if (1'b1) n467 <= 1'b0 ? 1'b0 : n855;
/* FF  7 12  1 */ always @(posedge clk) if (1'b1) n374 <= 1'b0 ? 1'b0 : n856;
/* FF  9 12  3 */ always @(posedge clk) if (1'b1) n513 <= 1'b0 ? 1'b0 : n857;
/* FF  5  4  4 */ assign n150 = n858;
/* FF  6  8  6 */ assign n264 = n859;
/* FF  7  4  6 */ assign n326 = n860;
/* FF  7 13  2 */ always @(posedge clk) if (1'b1) n382 <= 1'b0 ? 1'b0 : n861;
/* FF  5  5  5 */ assign n157 = n862;
/* FF  7  5  7 */ assign n169 = n863;
/* FF  8  4  1 */ assign n413 = n864;
/* FF  2  4  7 */ assign n59 = n865;
/* FF  6  7  1 */ assign n183 = n866;
/* FF  8  7  3 */ assign n435 = n867;
/* FF  5  8  6 */ always @(posedge clk) if (1'b1) n181 <= 1'b0 ? 1'b0 : n868;
/* FF  9  8  1 */ always @(posedge clk) if (1'b1) n493 <= 1'b0 ? 1'b0 : n869;
/* FF  5 11  2 */ always @(posedge clk) if (1'b1) n202 <= 1'b0 ? 1'b0 : n870;
/* FF  4  4  5 */ always @(posedge clk) if (1'b1) n107 <= 1'b0 ? 1'b0 : n871;
/* FF  7 11  4 */ always @(posedge clk) if (1'b1) n369 <= 1'b0 ? 1'b0 : n872;
/* FF  4  7  1 */ always @(posedge clk) if (1'b1) n117 <= 1'b0 ? 1'b0 : n873;
/* FF  1  3  4 */ always @(posedge clk) if (n53) n8 <= rst ? 1'b0 : n874;
/* FF  8 11  0 */ assign n463 = n875;
/* FF  6 11  7 */ always @(posedge clk) if (1'b1) n291 <= 1'b0 ? 1'b0 : n876;
/* FF 11  6  7 */ always @(posedge clk) if (1'b1) n536 <= 1'b0 ? 1'b0 : n877;
/* FF 11  9  3 */ always @(posedge clk) if (1'b1) n548 <= 1'b0 ? 1'b0 : n878;
/* FF  5 12  3 */ always @(posedge clk) if (1'b1) n210 <= 1'b0 ? 1'b0 : n879;
/* FF  7 12  5 */ always @(posedge clk) if (1'b1) n377 <= 1'b0 ? 1'b0 : n880;
/* FF  6  8  1 */ assign n260 = n881;
/* FF  4  8  2 */ always @(posedge clk) if (1'b1) n124 <= 1'b0 ? 1'b0 : n882;
/* FF  9 12  7 */ always @(posedge clk) if (1'b1) n517 <= 1'b0 ? 1'b0 : n883;
/* FF  8  8  3 */ assign n443 = n884;
/* FF  7  4  1 */ assign n323 = n885;
/* FF  5  5  0 */ assign n69 = n886;
/* FF  7  5  2 */ assign n330 = n887;
/* FF  9  5  4 */ always @(posedge clk) if (1'b1) n488 <= 1'b0 ? 1'b0 : n888;
/* FF  4 11  3 */ always @(posedge clk) if (1'b1) n140 <= 1'b0 ? 1'b0 : n889;
/* FF  2  3  6 */ assign n12 = n890;
/* FF  6  7  5 */ assign n257 = n891;
/* FF  8  7  7 */ assign n28 = n892;
/* FF  5  8  1 */ always @(posedge clk) if (1'b1) n177 <= 1'b0 ? 1'b0 : n893;
/* FF  7  8  3 */ assign n350 = n894;
/* FF  4  4  0 */ always @(posedge clk) if (1'b1) n105 <= 1'b0 ? 1'b0 : n895;
/* FF  9  8  5 */ always @(posedge clk) if (1'b1) n29 <= 1'b0 ? 1'b0 : n896;
/* FF  5 11  6 */ always @(posedge clk) if (1'b1) n205 <= 1'b0 ? 1'b0 : n897;
/* FF  4  7  5 */ always @(posedge clk) if (1'b1) n121 <= 1'b0 ? 1'b0 : n898;
/* FF  6 11  2 */ assign n286 = n899;
/* FF  8 11  4 */ always @(posedge clk) if (1'b1) n379 <= 1'b0 ? 1'b0 : n900;
/* FF 11  9  7 */ always @(posedge clk) if (1'b1) n506 <= 1'b0 ? 1'b0 : n901;
/* FF  7 12  0 */ always @(posedge clk) if (1'b1) n373 <= 1'b0 ? 1'b0 : n902;
/* FF  5 12  7 */ always @(posedge clk) if (1'b1) n213 <= 1'b0 ? 1'b0 : n903;
/* FF  9 12  2 */ always @(posedge clk) if (1'b1) n512 <= 1'b0 ? 1'b0 : n904;
/* FF  7  4  5 */ assign n325 = n905;
/* FF  8  3  5 */ assign n409 = n906;
/* FF  5  7  4 */ always @(posedge clk) if (1'b1) n162 <= n1 ? 1'b0 : n907;
/* FF  2  3  1 */ assign n51 = n908;
/* FF  4 11  7 */ always @(posedge clk) if (1'b1) n141 <= 1'b0 ? 1'b0 : n909;
/* FF  7  7  6 */ assign n347 = n910;
/* FF  4 14  3 */ always @(posedge clk) if (1'b1) n46 <= 1'b0 ? 1'b0 : n911;
/* FF  8  7  2 */ assign n176 = n912;
/* FF 11  5  5 */ always @(posedge clk) if (1'b1) n95 <= 1'b0 ? 1'b0 : n913;
/* FF  5  8  5 */ always @(posedge clk) if (1'b1) n180 <= 1'b0 ? 1'b0 : n914;
/* FF  9  8  0 */ always @(posedge clk) if (1'b1) n492 <= 1'b0 ? 1'b0 : n915;
/* FF  7  8  7 */ assign n352 = n916;
/* FF  5 11  1 */ always @(posedge clk) if (1'b1) n201 <= 1'b0 ? 1'b0 : n917;
/* FF  4  4  4 */ always @(posedge clk) if (1'b1) n106 <= 1'b0 ? 1'b0 : n918;
/* FF  7 11  3 */ always @(posedge clk) if (1'b1) n368 <= 1'b0 ? 1'b0 : n919;
/* FF  4  7  0 */ always @(posedge clk) if (1'b1) n116 <= 1'b0 ? 1'b0 : n920;
/* FF  1  3  3 */ always @(posedge clk) if (n53) n7 <= rst ? 1'b0 : n921;
/* FF  2  7  7 */ always @(posedge clk) if (1'b1) n70 <= n9 ? 1'b0 : n922;
/* FF 11  9  2 */ always @(posedge clk) if (1'b1) n547 <= 1'b0 ? 1'b0 : n923;
/* FF  5 12  2 */ always @(posedge clk) if (1'b1) n209 <= 1'b0 ? 1'b0 : n924;
/* FF  4  8  1 */ always @(posedge clk) if (1'b1) n123 <= 1'b0 ? 1'b0 : n925;
/* FF  9 12  6 */ always @(posedge clk) if (1'b1) n516 <= 1'b0 ? 1'b0 : n926;
/* FF  7  4  0 */ assign n322 = n927;
/* FF  2 11  4 */ always @(posedge clk) if (1'b1) n85 <= 1'b0 ? 1'b0 : n928;
/* FF 12 11  7 */ always @(posedge clk) if (1'b1) n86 <= 1'b0 ? 1'b0 : n929;
/* FF  8  3  0 */ assign n253 = n930;
/* FF  6  3  7 */ always @(posedge clk) if (n4) n231 <= 1'b0 ? 1'b0 : n931;
/* FF  4 11  2 */ always @(posedge clk) if (1'b1) n139 <= 1'b0 ? 1'b0 : n932;
/* FF  7  7  1 */ assign n343 = n933;
/* FF  2  3  5 */ assign n55 = n934;
/* FF  6  7  4 */ assign n27 = n935;
/* FF  8  7  6 */ assign n438 = n936;
/* FF  5  8  0 */ always @(posedge clk) if (1'b1) n172 <= 1'b0 ? 1'b0 : n937;
/* FF  7  8  2 */ assign n349 = n938;
/* FF 12 12  7 */ always @(posedge clk) if (1'b1) n532 <= n3 ? 1'b0 : n939;
/* FF  9  8  4 */ always @(posedge clk) if (1'b1) n496 <= 1'b0 ? 1'b0 : n940;
/* FF  5 11  5 */ always @(posedge clk) if (1'b1) n204 <= 1'b0 ? 1'b0 : n941;
/* FF  7 11  7 */ always @(posedge clk) if (1'b1) n214 <= 1'b0 ? 1'b0 : n942;
/* FF  4  7  4 */ always @(posedge clk) if (1'b1) n120 <= 1'b0 ? 1'b0 : n943;
/* FF 11  6  1 */ always @(posedge clk) if (1'b1) n535 <= 1'b0 ? 1'b0 : n944;
/* FF  5 14  7 */ always @(posedge clk) if (1'b1) n225 <= 1'b0 ? 1'b0 : n945;
/* FF  6 10  5 */ always @(posedge clk) if (1'b1) n282 <= 1'b0 ? 1'b0 : n946;
/* FF 11  9  6 */ always @(posedge clk) if (1'b1) n83 <= 1'b0 ? 1'b0 : n947;
/* FF  8 10  7 */ always @(posedge clk) if (1'b1) n460 <= 1'b0 ? 1'b0 : n948;
/* FF  6 13  1 */ always @(posedge clk) if (1'b1) n297 <= 1'b0 ? 1'b0 : n949;
/* FF  8  2  3 */ assign n401 = n950;
/* FF  9 11  5 */ always @(posedge clk) if (1'b1) n509 <= 1'b0 ? 1'b0 : n951;
/* FF 12 11  2 */ always @(posedge clk) if (1'b1) n557 <= 1'b0 ? 1'b0 : n952;
/* FF  5  6  2 */ assign \d_out[7]  = n953;
/* FF  4 10  5 */ always @(posedge clk) if (1'b1) n134 <= 1'b0 ? 1'b0 : n954;
/* FF  6  3  2 */ assign n229 = n955;
/* FF  8  3  4 */ assign n408 = n956;
/* FF 11 12  7 */ always @(posedge clk) if (1'b1) n41 <= 1'b0 ? 1'b0 : n957;
/* FF  2  3  0 */ assign n50 = n958;
/* FF  7  7  5 */ assign n346 = n959;
/* FF  4  3  2 */ always @(posedge clk) if (1'b1) n11 <= 1'b0 ? 1'b0 : n960;
/* FF  8  7  1 */ assign n434 = n961;
/* FF 11  5  4 */ always @(posedge clk) if (1'b1) n534 <= 1'b0 ? 1'b0 : n962;
/* FF  8  6  5 */ assign n429 = n963;
/* FF  5 11  0 */ assign n200 = n964;
/* FF  7 11  2 */ assign n367 = n965;
/* FF  2  6  1 */ assign n65 = n966;
/* FF  5 14  2 */ always @(posedge clk) if (1'b1) n223 <= 1'b0 ? 1'b0 : n967;
/* FF  6 10  0 */ always @(posedge clk) if (1'b1) n277 <= 1'b0 ? 1'b0 : n968;
/* FF  7 14  4 */ always @(posedge clk) if (1'b1) n392 <= 1'b0 ? 1'b0 : n969;
/* FF 11  9  1 */ always @(posedge clk) if (1'b1) n546 <= 1'b0 ? 1'b0 : n970;
/* FF  8 10  2 */ always @(posedge clk) if (1'b1) n455 <= 1'b0 ? 1'b0 : n971;
/* FF  9 14  6 */ always @(posedge clk) if (1'b1) n529 <= 1'b0 ? 1'b0 : n972;
/* FF  6 13  5 */ always @(posedge clk) if (1'b1) n301 <= 1'b0 ? 1'b0 : n973;
/* FF  8  2  7 */ assign n404 = n974;
/* FF  7  3  3 */ assign n319 = n975;
/* FF  4 10  0 */ always @(posedge clk) if (1'b1) n130 <= 1'b0 ? 1'b0 : n976;
/* FF  2 10  7 */ always @(posedge clk) if (1'b1) n82 <= 1'b0 ? 1'b0 : n977;
/* FF  5  6  6 */ always @(posedge clk) if (1'b1) n167 <= 1'b0 ? 1'b0 : n978;
/* FF  6 14  6 */ assign n3 = n979;
/* FF  6  3  6 */ assign n152 = n980;
/* FF  4  2  5 */ assign n103 = n981;
/* FF  6  6  2 */ always @(posedge clk) if (n4) n251 <= 1'b0 ? 1'b0 : n982;
/* FF  7 15  4 */ always @(posedge clk) if (1'b1) n396 <= 1'b0 ? 1'b0 : n983;
/* FF  4 11  1 */ always @(posedge clk) if (1'b1) n99 <= 1'b0 ? 1'b0 : n984;
/* FF  7  7  0 */ assign n342 = n985;
/* FF  2  3  4 */ assign n54 = n986;
/* FF  8  6  0 */ assign n425 = n987;
/* FF  6  9  3 */ assign n268 = n988;
/* FF  8  9  5 */ always @(posedge clk) if (1'b1) n450 <= 1'b0 ? 1'b0 : n989;
/* FF  2  6  5 */ assign n67 = n990;
/* FF  5 14  6 */ always @(posedge clk) if (1'b1) n224 <= 1'b0 ? 1'b0 : n991;
/* FF  9 14  1 */ always @(posedge clk) if (1'b1) n525 <= 1'b0 ? 1'b0 : n992;
/* FF  4  6  7 */ always @(posedge clk) if (1'b1) n113 <= n1 ? 1'b0 : n993;
/* FF  6 10  4 */ always @(posedge clk) if (1'b1) n281 <= 1'b0 ? 1'b0 : n994;
/* FF  8 10  6 */ always @(posedge clk) if (1'b1) n459 <= 1'b0 ? 1'b0 : n995;
/* FF  6 13  0 */ always @(posedge clk) if (1'b1) n296 <= 1'b0 ? 1'b0 : n996;
/* FF 11  8  0 */ assign \d_out[1]  = n997;
/* FF  8  2  2 */ assign n400 = n998;
/* FF  2 10  2 */ always @(posedge clk) if (1'b1) n79 <= 1'b0 ? 1'b0 : n999;
/* FF  7  3  7 */ assign n313 = n1000;
/* FF  4 10  4 */ always @(posedge clk) if (1'b1) n133 <= 1'b0 ? 1'b0 : n1001;
/* FF  8 14  3 */ always @(posedge clk) if (1'b1) n486 <= n3 ? 1'b0 : n1002;
/* FF 11 12  6 */ always @(posedge clk) if (1'b1) n87 <= 1'b0 ? 1'b0 : n1003;
/* FF  8 13  7 */ always @(posedge clk) if (1'b1) n484 <= 1'b0 ? 1'b0 : n1004;
/* FF  7  7  4 */ assign n345 = n1005;
/* FF  5 10  4 */ always @(posedge clk) if (1'b1) n197 <= 1'b0 ? 1'b0 : n1006;
/* FF  5 13  0 */ assign n215 = n1007;
/* FF  7 10  6 */ always @(posedge clk) if (1'b1) n39 <= 1'b0 ? 1'b0 : n1008;
/* FF  8  6  4 */ assign n428 = n1009;
/* FF  7  2  2 */ assign n306 = n1010;
/* FF  8  9  0 */ assign n446 = n1011;
/* FF  1  5  2 */ always @(posedge clk) if (1'b1) n13 <= n5 ? 1'b0 : n1012;
/* FF  6  9  7 */ always @(posedge clk) if (1'b1) n272 <= 1'b0 ? 1'b0 : n1013;
/* FF  2  6  0 */ assign n64 = n1014;
/* FF  5 14  1 */ always @(posedge clk) if (1'b1) n222 <= 1'b0 ? 1'b0 : n1015;
/* FF  4  6  2 */ assign n110 = n1016;
/* FF  7 14  3 */ always @(posedge clk) if (1'b1) n391 <= 1'b0 ? 1'b0 : n1017;
/* FF  8 10  1 */ always @(posedge clk) if (1'b1) n454 <= 1'b0 ? 1'b0 : n1018;
/* FF  9 14  5 */ always @(posedge clk) if (1'b1) n528 <= 1'b0 ? 1'b0 : n1019;
/* FF  6 13  4 */ always @(posedge clk) if (1'b1) n300 <= 1'b0 ? 1'b0 : n1020;
/* FF  8  2  6 */ assign n403 = n1021;
/* FF 11  8  4 */ always @(posedge clk) if (1'b1) n340 <= 1'b0 ? 1'b0 : n1022;
/* FF  7  3  2 */ assign n318 = n1023;
/* FF  2 10  6 */ always @(posedge clk) if (1'b1) n81 <= 1'b0 ? 1'b0 : n1024;
/* FF  5  6  5 */ always @(posedge clk) if (1'b1) n166 <= 1'b0 ? 1'b0 : n1025;
/* FF 12 11  5 */ always @(posedge clk) if (1'b1) n558 <= 1'b0 ? 1'b0 : n1026;
/* FF  2  2  2 */ always @(posedge clk) if (1'b1) n49 <= 1'b0 ? 1'b0 : n1027;
/* FF  7  6  4 */ assign n336 = n1028;
/* FF 11 12  1 */ always @(posedge clk) if (1'b1) n387 <= 1'b0 ? 1'b0 : n1029;
/* FF  8 13  2 */ always @(posedge clk) if (1'b1) n480 <= 1'b0 ? 1'b0 : n1030;
/* FF  5  9  7 */ always @(posedge clk) if (1'b1) n191 <= 1'b0 ? 1'b0 : n1031;
/* FF  2  5  4 */ always @(posedge clk) if (1'b1) n63 <= n5 ? 1'b0 : n1032;
/* FF  6  5  5 */ assign n246 = n1033;
/* FF  8  5  7 */ assign n424 = n1034;
/* FF  7 10  1 */ assign n360 = n1035;
/* FF  5 13  4 */ always @(posedge clk) if (1'b1) n219 <= 1'b0 ? 1'b0 : n1036;
/* FF  6  9  2 */ assign n267 = n1037;
/* FF  7  2  6 */ assign n310 = n1038;
/* FF  4  9  3 */ always @(posedge clk) if (1'b1) n36 <= 1'b0 ? 1'b0 : n1039;
/* FF  8  9  4 */ always @(posedge clk) if (1'b1) n449 <= 1'b0 ? 1'b0 : n1040;
/* FF 11  7  7 */ always @(posedge clk) if (1'b1) n541 <= 1'b0 ? 1'b0 : n1041;
/* FF  4  6  6 */ assign \d_out[6]  = n1042;
/* FF  8  2  1 */ assign n399 = n1043;
/* FF  6 12  3 */ assign n293 = n1044;
/* FF  8 12  5 */ always @(posedge clk) if (1'b1) n475 <= 1'b0 ? 1'b0 : n1045;
/* FF  5  6  0 */ assign n163 = n1046;
/* FF  5  9  2 */ always @(posedge clk) if (1'b1) n187 <= 1'b0 ? 1'b0 : n1047;
/* FF  6  5  0 */ assign n241 = n1048;
/* FF  8 13  6 */ always @(posedge clk) if (1'b1) n483 <= 1'b0 ? 1'b0 : n1049;
/* FF  4  5  1 */ always @(posedge clk) if (1'b1) n20 <= n5 ? 1'b0 : n1050;
/* FF  9  9  6 */ always @(posedge clk) if (1'b1) n502 <= 1'b0 ? 1'b0 : n1051;
/* FF  7  9  4 */ always @(posedge clk) if (1'b1) n356 <= 1'b0 ? 1'b0 : n1052;
/* FF  8  5  2 */ assign n419 = n1053;
/* FF 11  3  5 */ always @(posedge clk) if (1'b1) n487 <= 1'b0 ? 1'b0 : n1054;
/* FF  5 10  3 */ always @(posedge clk) if (1'b1) n37 <= 1'b0 ? 1'b0 : n1055;
/* FF  7 10  5 */ always @(posedge clk) if (1'b1) n363 <= 1'b0 ? 1'b0 : n1056;
/* FF  8  6  3 */ assign n427 = n1057;
/* FF  7  2  1 */ assign n305 = n1058;
/* FF  6  9  6 */ always @(posedge clk) if (1'b1) n271 <= 1'b0 ? 1'b0 : n1059;
/* FF  4  9  7 */ always @(posedge clk) if (1'b1) n84 <= 1'b0 ? 1'b0 : n1060;
/* FF 11  7  2 */ always @(posedge clk) if (1'b1) n539 <= 1'b0 ? 1'b0 : n1061;
/* FF  5 14  0 */ always @(posedge clk) if (1'b1) n221 <= 1'b0 ? 1'b0 : n1062;
/* FF  4  6  1 */ assign n109 = n1063;
/* FF  7 14  2 */ always @(posedge clk) if (1'b1) n390 <= 1'b0 ? 1'b0 : n1064;
/* FF  9 14  4 */ always @(posedge clk) if (1'b1) n527 <= 1'b0 ? 1'b0 : n1065;
/* FF  7 13  6 */ always @(posedge clk) if (1'b1) n380 <= 1'b0 ? 1'b0 : n1066;
/* FF 11  8  3 */ always @(posedge clk) if (1'b1) n333 <= 1'b0 ? 1'b0 : n1067;
/* FF  8 12  0 */ assign n471 = n1068;
/* FF  6 12  7 */ always @(posedge clk) if (1'b1) n295 <= 1'b0 ? 1'b0 : n1069;
/* FF  6  4  3 */ assign n234 = n1070;
/* FF  8  4  5 */ assign n416 = n1071;
/* FF  7  6  3 */ assign n335 = n1072;
/* FF  8 13  1 */ always @(posedge clk) if (1'b1) n479 <= 1'b0 ? 1'b0 : n1073;
/* FF  5  9  6 */ always @(posedge clk) if (1'b1) n190 <= 1'b0 ? 1'b0 : n1074;
/* FF  9  9  1 */ assign n38 = n1075;
/* FF  2  5  3 */ always @(posedge clk) if (1'b1) n62 <= n5 ? 1'b0 : n1076;
/* FF  6  5  4 */ assign n245 = n1077;
/* FF 11 11  4 */ always @(posedge clk) if (1'b1) n146 <= n3 ? 1'b0 : n1078;
/* FF  8  5  6 */ assign n423 = n1079;
/* FF  7 10  0 */ assign n265 = n1080;
/* FF  5 10  7 */ always @(posedge clk) if (1'b1) n199 <= 1'b0 ? 1'b0 : n1081;
/* FF  5 13  3 */ always @(posedge clk) if (1'b1) n218 <= 1'b0 ? 1'b0 : n1082;
/* FF  2  9  0 */ always @(posedge clk) if (1'b1) n75 <= 1'b0 ? 1'b0 : n1083;
/* FF  7  2  5 */ assign n309 = n1084;
/* FF  4  9  2 */ always @(posedge clk) if (1'b1) n35 <= 1'b0 ? 1'b0 : n1085;
/* FF  8  9  3 */ always @(posedge clk) if (1'b1) n448 <= 1'b0 ? 1'b0 : n1086;
/* FF  6  8  5 */ assign n254 = n1087;
/* FF  8  8  7 */ assign n273 = n1088;
/* FF  9 13  3 */ always @(posedge clk) if (1'b1) n520 <= 1'b0 ? 1'b0 : n1089;
/* FF  5  5  4 */ assign n156 = n1090;
/* FF  6 12  2 */ assign n292 = n1091;
/* FF  7  5  6 */ assign n327 = n1092;
/* FF  8 12  4 */ always @(posedge clk) if (1'b1) n474 <= 1'b0 ? 1'b0 : n1093;
/* FF  8  4  0 */ assign n412 = n1094;
/* FF  6  4  7 */ assign n237 = n1095;
/* FF  7  6  7 */ always @(posedge clk) if (n4) n338 <= 1'b0 ? 1'b0 : n1096;
/* FF  5  9  1 */ always @(posedge clk) if (1'b1) n186 <= 1'b0 ? 1'b0 : n1097;
/* FF  7  9  3 */ always @(posedge clk) if (1'b1) n32 <= 1'b0 ? 1'b0 : n1098;
/* FF  4  5  0 */ assign n18 = n1099;
/* FF  9  9  5 */ always @(posedge clk) if (1'b1) n501 <= 1'b0 ? 1'b0 : n1100;
/* FF  2  5  7 */ always @(posedge clk) if (1'b1) n22 <= n5 ? 1'b0 : n1101;
/* FF  8  5  1 */ assign n115 = n1102;
/* FF  7  2  0 */ assign n304 = n1103;
/* FF 11  7  1 */ always @(posedge clk) if (1'b1) n538 <= 1'b0 ? 1'b0 : n1104;
/* FF  8  8  2 */ assign n442 = n1105;
/* FF  7 13  5 */ always @(posedge clk) if (1'b1) n385 <= 1'b0 ? 1'b0 : n1106;
/* FF  7  5  1 */ assign n329 = n1107;
/* FF  9 13  7 */ always @(posedge clk) if (1'b1) n522 <= 1'b0 ? 1'b0 : n1108;
/* FF  6 12  6 */ always @(posedge clk) if (1'b1) n42 <= 1'b0 ? 1'b0 : n1109;
/* FF  6  4  2 */ assign n233 = n1110;
/* FF  8  4  4 */ assign n415 = n1111;
/* FF  7  6  2 */ assign n334 = n1112;
/* FF  9  9  0 */ assign n372 = n1113;
/* FF  2  5  2 */ always @(posedge clk) if (1'b1) n61 <= n5 ? 1'b0 : n1114;
/* FF 11 11  3 */ assign n518 = n1115;
/* FF  6 11  1 */ assign n288 = n1116;
/* FF  8 11  3 */ always @(posedge clk) if (1'b1) n466 <= 1'b0 ? 1'b0 : n1117;

endmodule

