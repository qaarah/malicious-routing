									// Reading file 'aes_select.asc'..

module chip (input clk, output d_vld, input rst, input select, output \d_out[5] , output \d_out[6] , output \d_out[7] , output \d_out[2] , output \d_out[4] , output \d_out[3] , output \d_out[0] , output \d_out[1] );

wire n1;
// (0, 0, 'glb_netwk_0')
// (2, 5, 'lutff_global/s_r')
// (2, 6, 'lutff_global/s_r')
// (4, 1, 'neigh_op_tnr_3')
// (4, 1, 'sp4_r_v_b_19')
// (4, 2, 'neigh_op_rgt_3')
// (4, 2, 'sp4_r_v_b_6')
// (4, 3, 'neigh_op_bnr_3')
// (4, 6, 'lutff_global/s_r')
// (5, 0, 'span4_horz_r_3')
// (5, 0, 'span4_vert_19')
// (5, 1, 'neigh_op_top_3')
// (5, 1, 'sp4_v_b_19')
// (5, 2, 'lutff_3/out')
// (5, 2, 'sp4_v_b_6')
// (5, 3, 'neigh_op_bot_3')
// (6, 0, 'span4_horz_r_7')
// (6, 1, 'neigh_op_tnl_3')
// (6, 2, 'neigh_op_lft_3')
// (6, 3, 'neigh_op_bnl_3')
// (7, 0, 'fabout')
// (7, 0, 'local_g0_3')
// (7, 0, 'span4_horz_r_11')
// (8, 0, 'span4_horz_r_15')
// (9, 0, 'span4_horz_l_15')

wire n2;
// (0, 0, 'glb_netwk_2')
// (4, 2, 'glb2local_1')
// (4, 2, 'local_g0_5')
// (4, 2, 'lutff_2/in_3')
// (6, 5, 'lutff_global/s_r')
// (6, 7, 'lutff_global/s_r')
// (8, 5, 'lutff_global/s_r')
// (8, 6, 'sp4_r_v_b_40')
// (8, 7, 'neigh_op_tnr_0')
// (8, 7, 'sp4_r_v_b_29')
// (8, 8, 'neigh_op_rgt_0')
// (8, 8, 'sp4_r_v_b_16')
// (8, 9, 'neigh_op_bnr_0')
// (8, 9, 'sp4_r_v_b_5')
// (9, 5, 'sp4_v_t_40')
// (9, 6, 'sp4_v_b_40')
// (9, 7, 'neigh_op_top_0')
// (9, 7, 'sp4_v_b_29')
// (9, 8, 'lutff_0/out')
// (9, 8, 'lutff_global/s_r')
// (9, 8, 'sp4_v_b_16')
// (9, 9, 'neigh_op_bot_0')
// (9, 9, 'sp4_h_r_5')
// (9, 9, 'sp4_v_b_5')
// (9, 13, 'lutff_global/s_r')
// (10, 7, 'neigh_op_tnl_0')
// (10, 8, 'neigh_op_lft_0')
// (10, 9, 'neigh_op_bnl_0')
// (10, 9, 'sp4_h_r_16')
// (11, 4, 'lutff_global/s_r')
// (11, 9, 'sp4_h_r_29')
// (12, 9, 'sp4_h_r_40')
// (13, 9, 'fabout')
// (13, 9, 'local_g1_0')
// (13, 9, 'span4_horz_40')

wire clk;
// (0, 0, 'glb_netwk_3')
// (0, 5, 'span4_vert_t_14')
// (0, 6, 'span4_vert_b_14')
// (0, 7, 'span4_vert_b_10')
// (0, 8, 'io_1/D_IN_0')
// (0, 8, 'io_1/PAD')
// (0, 8, 'span4_vert_b_6')
// (0, 9, 'fabout')
// (0, 9, 'local_g1_2')
// (0, 9, 'span4_vert_b_2')
// (1, 7, 'neigh_op_tnl_2')
// (1, 7, 'neigh_op_tnl_6')
// (1, 8, 'lutff_global/clk')
// (1, 8, 'neigh_op_lft_2')
// (1, 8, 'neigh_op_lft_6')
// (1, 9, 'neigh_op_bnl_2')
// (1, 9, 'neigh_op_bnl_6')
// (2, 2, 'lutff_global/clk')
// (2, 4, 'lutff_global/clk')
// (2, 5, 'lutff_global/clk')
// (2, 6, 'lutff_global/clk')
// (2, 7, 'lutff_global/clk')
// (2, 8, 'lutff_global/clk')
// (2, 9, 'lutff_global/clk')
// (2, 10, 'lutff_global/clk')
// (2, 11, 'lutff_global/clk')
// (2, 12, 'lutff_global/clk')
// (2, 13, 'lutff_global/clk')
// (2, 14, 'lutff_global/clk')
// (4, 2, 'lutff_global/clk')
// (4, 3, 'lutff_global/clk')
// (4, 5, 'lutff_global/clk')
// (4, 6, 'lutff_global/clk')
// (4, 9, 'lutff_global/clk')
// (4, 10, 'lutff_global/clk')
// (4, 11, 'lutff_global/clk')
// (4, 12, 'lutff_global/clk')
// (4, 13, 'lutff_global/clk')
// (4, 14, 'lutff_global/clk')
// (5, 2, 'lutff_global/clk')
// (5, 5, 'lutff_global/clk')
// (5, 8, 'lutff_global/clk')
// (5, 9, 'lutff_global/clk')
// (5, 10, 'lutff_global/clk')
// (5, 11, 'lutff_global/clk')
// (5, 12, 'lutff_global/clk')
// (5, 13, 'lutff_global/clk')
// (5, 14, 'lutff_global/clk')
// (6, 5, 'lutff_global/clk')
// (6, 6, 'lutff_global/clk')
// (6, 7, 'lutff_global/clk')
// (6, 8, 'lutff_global/clk')
// (6, 9, 'lutff_global/clk')
// (6, 10, 'lutff_global/clk')
// (6, 11, 'lutff_global/clk')
// (6, 12, 'lutff_global/clk')
// (6, 13, 'lutff_global/clk')
// (6, 14, 'lutff_global/clk')
// (6, 15, 'lutff_global/clk')
// (7, 5, 'lutff_global/clk')
// (7, 6, 'lutff_global/clk')
// (7, 7, 'lutff_global/clk')
// (7, 8, 'lutff_global/clk')
// (7, 9, 'lutff_global/clk')
// (7, 10, 'lutff_global/clk')
// (7, 11, 'lutff_global/clk')
// (7, 12, 'lutff_global/clk')
// (7, 13, 'lutff_global/clk')
// (7, 14, 'lutff_global/clk')
// (7, 15, 'lutff_global/clk')
// (8, 5, 'lutff_global/clk')
// (8, 6, 'lutff_global/clk')
// (8, 7, 'lutff_global/clk')
// (8, 8, 'lutff_global/clk')
// (8, 9, 'lutff_global/clk')
// (8, 10, 'lutff_global/clk')
// (8, 11, 'lutff_global/clk')
// (8, 12, 'lutff_global/clk')
// (8, 13, 'lutff_global/clk')
// (9, 5, 'lutff_global/clk')
// (9, 6, 'lutff_global/clk')
// (9, 7, 'lutff_global/clk')
// (9, 8, 'lutff_global/clk')
// (9, 9, 'lutff_global/clk')
// (9, 10, 'lutff_global/clk')
// (9, 11, 'lutff_global/clk')
// (9, 12, 'lutff_global/clk')
// (9, 13, 'lutff_global/clk')
// (11, 4, 'lutff_global/clk')
// (11, 5, 'lutff_global/clk')
// (11, 6, 'lutff_global/clk')
// (11, 7, 'lutff_global/clk')
// (11, 8, 'lutff_global/clk')
// (11, 9, 'lutff_global/clk')
// (11, 10, 'lutff_global/clk')
// (11, 11, 'lutff_global/clk')
// (11, 12, 'lutff_global/clk')
// (11, 13, 'lutff_global/clk')
// (12, 6, 'lutff_global/clk')
// (12, 7, 'lutff_global/clk')
// (12, 9, 'lutff_global/clk')

reg n4 = 0;
// (0, 0, 'glb_netwk_5')
// (2, 2, 'glb2local_0')
// (2, 2, 'local_g0_4')
// (2, 2, 'lutff_4/in_2')
// (2, 4, 'glb2local_0')
// (2, 4, 'local_g0_4')
// (2, 4, 'lutff_1/in_3')
// (2, 4, 'lutff_global/cen')
// (4, 1, 'neigh_op_tnr_7')
// (4, 2, 'neigh_op_rgt_7')
// (4, 3, 'neigh_op_bnr_7')
// (5, 1, 'neigh_op_top_7')
// (5, 1, 'sp4_r_v_b_26')
// (5, 2, 'lutff_7/out')
// (5, 2, 'sp4_r_v_b_15')
// (5, 3, 'glb2local_1')
// (5, 3, 'local_g0_5')
// (5, 3, 'lutff_3/in_0')
// (5, 3, 'neigh_op_bot_7')
// (5, 3, 'sp4_r_v_b_2')
// (6, 0, 'fabout')
// (6, 0, 'local_g1_2')
// (6, 0, 'span4_vert_26')
// (6, 1, 'neigh_op_tnl_7')
// (6, 1, 'sp4_v_b_26')
// (6, 2, 'neigh_op_lft_7')
// (6, 2, 'sp4_v_b_15')
// (6, 3, 'neigh_op_bnl_7')
// (6, 3, 'sp4_v_b_2')
// (6, 4, 'glb2local_1')
// (6, 4, 'glb2local_2')
// (6, 4, 'local_g0_5')
// (6, 4, 'local_g0_6')
// (6, 4, 'lutff_2/in_3')
// (6, 4, 'lutff_5/in_3')
// (6, 5, 'glb2local_0')
// (6, 5, 'glb2local_3')
// (6, 5, 'local_g0_4')
// (6, 5, 'local_g0_7')
// (6, 5, 'lutff_2/in_3')
// (6, 5, 'lutff_3/in_3')
// (6, 5, 'lutff_4/in_3')
// (7, 5, 'glb2local_1')
// (7, 5, 'local_g0_5')
// (7, 5, 'lutff_0/in_3')
// (7, 6, 'lutff_global/cen')
// (9, 5, 'lutff_global/cen')
// (11, 6, 'lutff_global/cen')

wire n5;
// (0, 0, 'glb_netwk_6')
// (0, 8, 'fabout')
// (0, 8, 'local_g0_1')
// (0, 8, 'span4_horz_25')
// (1, 8, 'sp4_h_r_36')
// (2, 8, 'sp4_h_l_36')
// (2, 8, 'sp4_h_r_10')
// (2, 10, 'lutff_global/s_r')
// (3, 7, 'neigh_op_tnr_1')
// (3, 8, 'neigh_op_rgt_1')
// (3, 8, 'sp4_h_r_23')
// (3, 9, 'neigh_op_bnr_1')
// (4, 7, 'neigh_op_top_1')
// (4, 8, 'lutff_1/out')
// (4, 8, 'sp4_h_r_34')
// (4, 9, 'neigh_op_bot_1')
// (5, 7, 'neigh_op_tnl_1')
// (5, 8, 'lutff_global/s_r')
// (5, 8, 'neigh_op_lft_1')
// (5, 8, 'sp4_h_r_47')
// (5, 9, 'lutff_global/s_r')
// (5, 9, 'neigh_op_bnl_1')
// (5, 10, 'lutff_global/s_r')
// (6, 8, 'sp4_h_l_47')

reg n6 = 0;
// (0, 2, 'span12_horz_0')
// (1, 1, 'neigh_op_tnr_6')
// (1, 2, 'neigh_op_rgt_6')
// (1, 2, 'sp12_h_r_3')
// (1, 2, 'sp4_h_r_3')
// (1, 3, 'neigh_op_bnr_6')
// (2, 1, 'neigh_op_top_6')
// (2, 1, 'sp4_r_v_b_24')
// (2, 2, 'lutff_6/out')
// (2, 2, 'sp12_h_r_4')
// (2, 2, 'sp4_h_r_14')
// (2, 2, 'sp4_r_v_b_13')
// (2, 3, 'neigh_op_bot_6')
// (2, 3, 'sp4_r_v_b_0')
// (3, 0, 'span4_vert_24')
// (3, 1, 'neigh_op_tnl_6')
// (3, 1, 'sp4_v_b_24')
// (3, 2, 'neigh_op_lft_6')
// (3, 2, 'sp12_h_r_7')
// (3, 2, 'sp4_h_r_27')
// (3, 2, 'sp4_v_b_13')
// (3, 3, 'neigh_op_bnl_6')
// (3, 3, 'sp4_h_r_0')
// (3, 3, 'sp4_v_b_0')
// (4, 2, 'local_g1_0')
// (4, 2, 'lutff_7/in_2')
// (4, 2, 'sp12_h_r_8')
// (4, 2, 'sp4_h_r_38')
// (4, 3, 'sp4_h_r_13')
// (4, 3, 'sp4_r_v_b_45')
// (4, 4, 'sp4_r_v_b_32')
// (4, 5, 'sp4_r_v_b_21')
// (4, 6, 'sp4_r_v_b_8')
// (5, 2, 'sp12_h_r_11')
// (5, 2, 'sp4_h_l_38')
// (5, 2, 'sp4_h_r_0')
// (5, 2, 'sp4_h_r_1')
// (5, 2, 'sp4_v_t_45')
// (5, 3, 'local_g2_0')
// (5, 3, 'lutff_3/in_1')
// (5, 3, 'sp4_h_r_24')
// (5, 3, 'sp4_v_b_45')
// (5, 4, 'local_g2_0')
// (5, 4, 'lutff_1/in_1')
// (5, 4, 'sp4_v_b_32')
// (5, 5, 'sp4_v_b_21')
// (5, 6, 'sp4_v_b_8')
// (6, 2, 'sp12_h_r_12')
// (6, 2, 'sp4_h_r_12')
// (6, 2, 'sp4_h_r_13')
// (6, 3, 'sp4_h_r_37')
// (6, 4, 'sp4_r_v_b_40')
// (6, 5, 'sp4_r_v_b_29')
// (6, 6, 'sp4_r_v_b_16')
// (6, 7, 'sp4_r_v_b_5')
// (7, 2, 'sp12_h_r_15')
// (7, 2, 'sp4_h_r_24')
// (7, 2, 'sp4_h_r_25')
// (7, 3, 'sp4_h_l_37')
// (7, 3, 'sp4_h_r_8')
// (7, 3, 'sp4_v_t_40')
// (7, 4, 'local_g2_0')
// (7, 4, 'lutff_7/in_1')
// (7, 4, 'sp4_v_b_40')
// (7, 5, 'local_g2_5')
// (7, 5, 'lutff_4/in_1')
// (7, 5, 'sp4_v_b_29')
// (7, 6, 'sp4_v_b_16')
// (7, 7, 'sp4_v_b_5')
// (8, 2, 'sp12_h_r_16')
// (8, 2, 'sp4_h_r_36')
// (8, 2, 'sp4_h_r_37')
// (8, 3, 'sp4_h_r_21')
// (8, 3, 'sp4_r_v_b_36')
// (8, 3, 'sp4_r_v_b_37')
// (8, 3, 'sp4_r_v_b_43')
// (8, 4, 'sp4_r_v_b_24')
// (8, 4, 'sp4_r_v_b_25')
// (8, 4, 'sp4_r_v_b_30')
// (8, 5, 'local_g2_4')
// (8, 5, 'local_g2_5')
// (8, 5, 'lutff_1/in_1')
// (8, 5, 'lutff_4/in_1')
// (8, 5, 'lutff_6/in_1')
// (8, 5, 'sp4_r_v_b_12')
// (8, 5, 'sp4_r_v_b_13')
// (8, 5, 'sp4_r_v_b_19')
// (8, 6, 'sp4_r_v_b_0')
// (8, 6, 'sp4_r_v_b_1')
// (8, 6, 'sp4_r_v_b_6')
// (9, 2, 'sp12_h_r_19')
// (9, 2, 'sp4_h_l_36')
// (9, 2, 'sp4_h_l_37')
// (9, 2, 'sp4_v_t_36')
// (9, 2, 'sp4_v_t_37')
// (9, 2, 'sp4_v_t_43')
// (9, 3, 'sp4_h_r_32')
// (9, 3, 'sp4_v_b_36')
// (9, 3, 'sp4_v_b_37')
// (9, 3, 'sp4_v_b_43')
// (9, 4, 'local_g3_1')
// (9, 4, 'lutff_5/in_1')
// (9, 4, 'sp4_v_b_24')
// (9, 4, 'sp4_v_b_25')
// (9, 4, 'sp4_v_b_30')
// (9, 5, 'local_g1_3')
// (9, 5, 'local_g1_4')
// (9, 5, 'lutff_1/in_2')
// (9, 5, 'lutff_4/in_1')
// (9, 5, 'lutff_5/in_1')
// (9, 5, 'sp4_v_b_12')
// (9, 5, 'sp4_v_b_13')
// (9, 5, 'sp4_v_b_19')
// (9, 6, 'sp4_v_b_0')
// (9, 6, 'sp4_v_b_1')
// (9, 6, 'sp4_v_b_6')
// (10, 2, 'sp12_h_r_20')
// (10, 3, 'sp4_h_r_45')
// (10, 4, 'sp4_r_v_b_36')
// (10, 5, 'sp4_r_v_b_25')
// (10, 6, 'sp4_r_v_b_12')
// (10, 7, 'sp4_r_v_b_1')
// (11, 2, 'sp12_h_r_23')
// (11, 3, 'sp4_h_l_45')
// (11, 3, 'sp4_r_v_b_45')
// (11, 3, 'sp4_v_t_36')
// (11, 4, 'local_g0_3')
// (11, 4, 'lutff_2/in_1')
// (11, 4, 'lutff_6/in_1')
// (11, 4, 'sp4_r_v_b_32')
// (11, 4, 'sp4_v_b_36')
// (11, 5, 'local_g2_1')
// (11, 5, 'local_g3_5')
// (11, 5, 'lutff_0/in_1')
// (11, 5, 'lutff_1/in_1')
// (11, 5, 'lutff_3/in_1')
// (11, 5, 'sp4_r_v_b_21')
// (11, 5, 'sp4_v_b_25')
// (11, 6, 'sp4_r_v_b_8')
// (11, 6, 'sp4_v_b_12')
// (11, 7, 'sp4_v_b_1')
// (12, 2, 'sp12_h_l_23')
// (12, 2, 'sp12_v_t_23')
// (12, 2, 'sp4_v_t_45')
// (12, 3, 'sp12_v_b_23')
// (12, 3, 'sp4_v_b_45')
// (12, 4, 'sp12_v_b_20')
// (12, 4, 'sp4_v_b_32')
// (12, 5, 'sp12_v_b_19')
// (12, 5, 'sp4_v_b_21')
// (12, 6, 'sp12_v_b_16')
// (12, 6, 'sp4_v_b_8')
// (12, 7, 'sp12_v_b_15')
// (12, 8, 'sp12_v_b_12')
// (12, 9, 'sp12_v_b_11')
// (12, 10, 'sp12_v_b_8')
// (12, 11, 'sp12_v_b_7')
// (12, 12, 'sp12_v_b_4')
// (12, 13, 'sp12_v_b_3')
// (12, 14, 'sp12_v_b_0')

wire n7;
// (0, 2, 'span12_horz_10')
// (1, 2, 'sp12_h_r_13')
// (2, 2, 'sp12_h_r_14')
// (3, 2, 'sp12_h_r_17')
// (4, 2, 'sp12_h_r_18')
// (4, 3, 'sp4_r_v_b_47')
// (4, 4, 'sp4_r_v_b_34')
// (4, 5, 'sp4_r_v_b_23')
// (4, 6, 'sp4_r_v_b_10')
// (4, 7, 'sp4_r_v_b_47')
// (4, 8, 'sp4_r_v_b_34')
// (4, 9, 'sp4_r_v_b_23')
// (4, 10, 'sp4_r_v_b_10')
// (5, 2, 'sp12_h_r_21')
// (5, 2, 'sp4_h_r_10')
// (5, 2, 'sp4_v_t_47')
// (5, 3, 'sp4_v_b_47')
// (5, 4, 'sp4_v_b_34')
// (5, 5, 'sp4_v_b_23')
// (5, 6, 'local_g0_2')
// (5, 6, 'lutff_1/in_1')
// (5, 6, 'lutff_2/in_2')
// (5, 6, 'sp4_v_b_10')
// (5, 6, 'sp4_v_t_47')
// (5, 7, 'sp4_v_b_47')
// (5, 8, 'local_g2_2')
// (5, 8, 'lutff_1/in_3')
// (5, 8, 'sp4_v_b_34')
// (5, 9, 'sp4_v_b_23')
// (5, 10, 'sp4_v_b_10')
// (6, 2, 'sp12_h_r_22')
// (6, 2, 'sp4_h_r_23')
// (6, 6, 'sp4_r_v_b_42')
// (6, 7, 'local_g1_7')
// (6, 7, 'lutff_2/in_2')
// (6, 7, 'sp4_r_v_b_31')
// (6, 8, 'sp4_r_v_b_18')
// (6, 9, 'sp4_r_v_b_7')
// (6, 12, 'neigh_op_tnr_1')
// (6, 13, 'neigh_op_rgt_1')
// (6, 14, 'neigh_op_bnr_1')
// (7, 2, 'sp12_h_l_22')
// (7, 2, 'sp12_v_t_22')
// (7, 2, 'sp4_h_r_34')
// (7, 3, 'sp12_v_b_22')
// (7, 4, 'sp12_v_b_21')
// (7, 5, 'sp12_v_b_18')
// (7, 5, 'sp4_v_t_42')
// (7, 6, 'sp12_v_b_17')
// (7, 6, 'sp4_v_b_42')
// (7, 7, 'sp12_v_b_14')
// (7, 7, 'sp4_v_b_31')
// (7, 8, 'sp12_v_b_13')
// (7, 8, 'sp4_v_b_18')
// (7, 9, 'local_g3_2')
// (7, 9, 'lutff_3/in_2')
// (7, 9, 'sp12_v_b_10')
// (7, 9, 'sp4_v_b_7')
// (7, 10, 'sp12_v_b_9')
// (7, 11, 'sp12_v_b_6')
// (7, 12, 'neigh_op_top_1')
// (7, 12, 'sp12_v_b_5')
// (7, 13, 'lutff_1/out')
// (7, 13, 'sp12_v_b_2')
// (7, 14, 'neigh_op_bot_1')
// (7, 14, 'sp12_v_b_1')
// (8, 2, 'sp4_h_r_47')
// (8, 12, 'neigh_op_tnl_1')
// (8, 13, 'neigh_op_lft_1')
// (8, 14, 'neigh_op_bnl_1')
// (9, 2, 'sp4_h_l_47')

reg n8 = 0;
// (0, 2, 'span4_horz_0')
// (1, 1, 'neigh_op_tnr_4')
// (1, 2, 'neigh_op_rgt_4')
// (1, 2, 'sp4_h_r_13')
// (1, 3, 'neigh_op_bnr_4')
// (2, 1, 'neigh_op_top_4')
// (2, 2, 'local_g1_4')
// (2, 2, 'lutff_4/in_1')
// (2, 2, 'lutff_4/out')
// (2, 2, 'lutff_6/in_3')
// (2, 2, 'sp4_h_r_24')
// (2, 2, 'sp4_h_r_8')
// (2, 3, 'neigh_op_bot_4')
// (3, 1, 'neigh_op_tnl_4')
// (3, 2, 'neigh_op_lft_4')
// (3, 2, 'sp4_h_r_21')
// (3, 2, 'sp4_h_r_37')
// (3, 3, 'neigh_op_bnl_4')
// (3, 3, 'sp4_r_v_b_40')
// (3, 4, 'sp4_r_v_b_29')
// (3, 5, 'sp4_r_v_b_16')
// (3, 6, 'sp4_r_v_b_5')
// (4, 2, 'local_g2_0')
// (4, 2, 'lutff_1/in_1')
// (4, 2, 'sp4_h_l_37')
// (4, 2, 'sp4_h_r_32')
// (4, 2, 'sp4_v_t_40')
// (4, 3, 'local_g2_0')
// (4, 3, 'lutff_4/in_0')
// (4, 3, 'sp4_v_b_40')
// (4, 4, 'sp4_v_b_29')
// (4, 5, 'sp4_v_b_16')
// (4, 6, 'sp4_v_b_5')
// (5, 2, 'sp4_h_r_45')
// (5, 3, 'local_g2_4')
// (5, 3, 'lutff_3/in_3')
// (5, 3, 'sp4_r_v_b_36')
// (5, 4, 'sp4_r_v_b_25')
// (5, 5, 'sp4_r_v_b_12')
// (5, 6, 'sp4_r_v_b_1')
// (6, 2, 'sp4_h_l_45')
// (6, 2, 'sp4_v_t_36')
// (6, 3, 'sp4_v_b_36')
// (6, 4, 'sp4_v_b_25')
// (6, 5, 'sp4_v_b_12')
// (6, 6, 'sp4_v_b_1')

wire n9;
// (0, 3, 'span12_horz_6')
// (1, 3, 'sp12_h_r_9')
// (2, 3, 'sp12_h_r_10')
// (3, 3, 'sp12_h_r_13')
// (4, 3, 'sp12_h_r_14')
// (5, 2, 'neigh_op_tnr_5')
// (5, 3, 'neigh_op_rgt_5')
// (5, 3, 'sp12_h_r_17')
// (5, 4, 'neigh_op_bnr_5')
// (6, 2, 'neigh_op_top_5')
// (6, 3, 'lutff_5/out')
// (6, 3, 'sp12_h_r_18')
// (6, 4, 'neigh_op_bot_5')
// (7, 2, 'neigh_op_tnl_5')
// (7, 3, 'neigh_op_lft_5')
// (7, 3, 'sp12_h_r_21')
// (7, 3, 'sp4_h_r_10')
// (7, 4, 'local_g2_5')
// (7, 4, 'local_g3_5')
// (7, 4, 'lutff_0/in_2')
// (7, 4, 'lutff_5/in_2')
// (7, 4, 'neigh_op_bnl_5')
// (8, 3, 'local_g0_6')
// (8, 3, 'local_g0_7')
// (8, 3, 'lutff_0/in_2')
// (8, 3, 'lutff_6/in_3')
// (8, 3, 'sp12_h_r_22')
// (8, 3, 'sp4_h_r_23')
// (9, 3, 'sp12_h_l_22')
// (9, 3, 'sp4_h_r_34')
// (10, 3, 'sp4_h_r_47')
// (11, 3, 'sp4_h_l_47')

wire n10;
// (0, 4, 'span12_horz_1')
// (1, 4, 'sp12_h_r_2')
// (2, 4, 'sp12_h_r_5')
// (3, 4, 'sp12_h_r_6')
// (4, 4, 'sp12_h_r_9')
// (5, 4, 'sp12_h_r_10')
// (6, 3, 'neigh_op_tnr_3')
// (6, 4, 'neigh_op_rgt_3')
// (6, 4, 'sp12_h_r_13')
// (6, 5, 'neigh_op_bnr_3')
// (7, 3, 'neigh_op_top_3')
// (7, 4, 'lutff_3/out')
// (7, 4, 'sp12_h_r_14')
// (7, 5, 'neigh_op_bot_3')
// (8, 3, 'neigh_op_tnl_3')
// (8, 4, 'local_g0_1')
// (8, 4, 'lutff_7/in_2')
// (8, 4, 'neigh_op_lft_3')
// (8, 4, 'sp12_h_r_17')
// (8, 5, 'neigh_op_bnl_3')
// (9, 4, 'sp12_h_r_18')
// (10, 4, 'sp12_h_r_21')
// (11, 4, 'sp12_h_r_22')
// (12, 4, 'sp12_h_l_22')

reg n11 = 0;
// (0, 4, 'span12_horz_12')
// (1, 3, 'neigh_op_tnr_4')
// (1, 4, 'neigh_op_rgt_4')
// (1, 4, 'sp12_h_r_15')
// (1, 5, 'neigh_op_bnr_4')
// (2, 3, 'neigh_op_top_4')
// (2, 4, 'lutff_4/out')
// (2, 4, 'sp12_h_r_16')
// (2, 5, 'neigh_op_bot_4')
// (3, 3, 'neigh_op_tnl_4')
// (3, 4, 'neigh_op_lft_4')
// (3, 4, 'sp12_h_r_19')
// (3, 5, 'neigh_op_bnl_4')
// (4, 4, 'sp12_h_r_20')
// (5, 4, 'local_g1_7')
// (5, 4, 'lutff_1/in_3')
// (5, 4, 'sp12_h_r_23')
// (6, 4, 'sp12_h_l_23')

wire n12;
// (0, 4, 'span12_horz_2')
// (1, 4, 'sp12_h_r_5')
// (2, 4, 'sp12_h_r_6')
// (3, 4, 'sp12_h_r_9')
// (4, 4, 'sp12_h_r_10')
// (4, 5, 'sp12_h_r_1')
// (5, 4, 'sp12_h_r_13')
// (5, 5, 'sp12_h_r_2')
// (6, 4, 'sp12_h_r_14')
// (6, 5, 'sp12_h_r_5')
// (7, 4, 'sp12_h_r_17')
// (7, 5, 'sp12_h_r_6')
// (8, 4, 'sp12_h_r_18')
// (8, 5, 'sp12_h_r_9')
// (9, 4, 'local_g0_5')
// (9, 4, 'lutff_3/in_2')
// (9, 4, 'sp12_h_r_21')
// (9, 5, 'local_g1_2')
// (9, 5, 'lutff_3/in_2')
// (9, 5, 'sp12_h_r_10')
// (10, 4, 'neigh_op_tnr_3')
// (10, 4, 'sp12_h_r_22')
// (10, 5, 'neigh_op_rgt_3')
// (10, 5, 'sp12_h_r_13')
// (10, 6, 'neigh_op_bnr_3')
// (11, 4, 'neigh_op_top_3')
// (11, 4, 'sp12_h_l_22')
// (11, 4, 'sp12_v_t_22')
// (11, 5, 'lutff_3/out')
// (11, 5, 'sp12_h_r_14')
// (11, 5, 'sp12_v_b_22')
// (11, 6, 'neigh_op_bot_3')
// (11, 6, 'sp12_v_b_21')
// (11, 7, 'sp12_v_b_18')
// (11, 8, 'sp12_v_b_17')
// (11, 9, 'sp12_v_b_14')
// (11, 10, 'sp12_v_b_13')
// (11, 11, 'sp12_v_b_10')
// (11, 12, 'sp12_v_b_9')
// (11, 13, 'sp12_v_b_6')
// (11, 14, 'sp12_v_b_5')
// (11, 15, 'sp12_v_b_2')
// (11, 16, 'sp12_v_b_1')
// (12, 4, 'neigh_op_tnl_3')
// (12, 5, 'neigh_op_lft_3')
// (12, 5, 'sp12_h_r_17')
// (12, 6, 'neigh_op_bnl_3')
// (13, 5, 'span12_horz_17')

wire n13;
// (0, 4, 'span12_horz_6')
// (1, 4, 'sp12_h_r_9')
// (2, 4, 'sp12_h_r_10')
// (3, 4, 'sp12_h_r_13')
// (4, 4, 'sp12_h_r_14')
// (5, 3, 'neigh_op_tnr_5')
// (5, 4, 'neigh_op_rgt_5')
// (5, 4, 'sp12_h_r_17')
// (5, 5, 'neigh_op_bnr_5')
// (6, 3, 'neigh_op_top_5')
// (6, 4, 'local_g1_2')
// (6, 4, 'lutff_0/in_3')
// (6, 4, 'lutff_5/out')
// (6, 4, 'lutff_6/in_3')
// (6, 4, 'sp12_h_r_18')
// (6, 5, 'neigh_op_bot_5')
// (7, 3, 'neigh_op_tnl_5')
// (7, 4, 'neigh_op_lft_5')
// (7, 4, 'sp12_h_r_21')
// (7, 5, 'neigh_op_bnl_5')
// (8, 4, 'sp12_h_r_22')
// (9, 4, 'sp12_h_l_22')

reg n14 = 0;
// (0, 5, 'span12_horz_2')
// (1, 4, 'neigh_op_tnr_7')
// (1, 5, 'neigh_op_rgt_7')
// (1, 5, 'sp12_h_r_5')
// (1, 6, 'neigh_op_bnr_7')
// (2, 4, 'local_g1_7')
// (2, 4, 'lutff_2/in_2')
// (2, 4, 'lutff_3/in_1')
// (2, 4, 'neigh_op_top_7')
// (2, 5, 'local_g2_7')
// (2, 5, 'lutff_7/in_2')
// (2, 5, 'lutff_7/out')
// (2, 5, 'sp12_h_r_6')
// (2, 6, 'neigh_op_bot_7')
// (3, 4, 'neigh_op_tnl_7')
// (3, 5, 'neigh_op_lft_7')
// (3, 5, 'sp12_h_r_9')
// (3, 5, 'sp4_h_r_4')
// (3, 6, 'neigh_op_bnl_7')
// (4, 2, 'sp4_r_v_b_43')
// (4, 3, 'sp4_r_v_b_30')
// (4, 4, 'sp4_r_v_b_19')
// (4, 5, 'sp12_h_r_10')
// (4, 5, 'sp4_h_r_17')
// (4, 5, 'sp4_r_v_b_6')
// (5, 1, 'sp4_v_t_43')
// (5, 2, 'sp4_v_b_43')
// (5, 3, 'sp4_v_b_30')
// (5, 4, 'local_g0_3')
// (5, 4, 'lutff_5/in_2')
// (5, 4, 'sp4_v_b_19')
// (5, 5, 'sp12_h_r_13')
// (5, 5, 'sp4_h_r_28')
// (5, 5, 'sp4_h_r_6')
// (5, 5, 'sp4_v_b_6')
// (6, 1, 'sp4_r_v_b_4')
// (6, 2, 'sp4_r_v_b_41')
// (6, 2, 'sp4_r_v_b_42')
// (6, 3, 'sp4_r_v_b_28')
// (6, 3, 'sp4_r_v_b_31')
// (6, 4, 'local_g3_1')
// (6, 4, 'local_g3_2')
// (6, 4, 'lutff_0/in_0')
// (6, 4, 'lutff_2/in_0')
// (6, 4, 'lutff_5/in_2')
// (6, 4, 'sp4_r_v_b_17')
// (6, 4, 'sp4_r_v_b_18')
// (6, 5, 'local_g1_3')
// (6, 5, 'local_g1_6')
// (6, 5, 'lutff_3/in_1')
// (6, 5, 'lutff_5/in_2')
// (6, 5, 'lutff_6/in_2')
// (6, 5, 'sp12_h_r_14')
// (6, 5, 'sp4_h_r_19')
// (6, 5, 'sp4_h_r_41')
// (6, 5, 'sp4_r_v_b_4')
// (6, 5, 'sp4_r_v_b_7')
// (7, 0, 'span4_vert_4')
// (7, 1, 'sp4_v_b_4')
// (7, 1, 'sp4_v_t_41')
// (7, 1, 'sp4_v_t_42')
// (7, 2, 'sp4_v_b_41')
// (7, 2, 'sp4_v_b_42')
// (7, 3, 'sp4_v_b_28')
// (7, 3, 'sp4_v_b_31')
// (7, 4, 'sp4_v_b_17')
// (7, 4, 'sp4_v_b_18')
// (7, 5, 'sp12_h_r_17')
// (7, 5, 'sp4_h_l_41')
// (7, 5, 'sp4_h_r_30')
// (7, 5, 'sp4_v_b_4')
// (7, 5, 'sp4_v_b_7')
// (8, 5, 'sp12_h_r_18')
// (8, 5, 'sp4_h_r_43')
// (9, 5, 'sp12_h_r_21')
// (9, 5, 'sp4_h_l_43')
// (10, 5, 'sp12_h_r_22')
// (11, 5, 'sp12_h_l_22')

reg n15 = 0;
// (0, 5, 'span12_horz_7')
// (1, 5, 'sp12_h_r_8')
// (2, 5, 'sp12_h_r_11')
// (3, 5, 'sp12_h_r_12')
// (4, 4, 'neigh_op_tnr_4')
// (4, 5, 'neigh_op_rgt_4')
// (4, 5, 'sp12_h_r_15')
// (4, 6, 'neigh_op_bnr_4')
// (5, 4, 'neigh_op_top_4')
// (5, 5, 'lutff_4/out')
// (5, 5, 'sp12_h_r_16')
// (5, 5, 'sp4_h_r_8')
// (5, 6, 'neigh_op_bot_4')
// (6, 4, 'neigh_op_tnl_4')
// (6, 5, 'neigh_op_lft_4')
// (6, 5, 'sp12_h_r_19')
// (6, 5, 'sp4_h_r_21')
// (6, 6, 'neigh_op_bnl_4')
// (7, 5, 'sp12_h_r_20')
// (7, 5, 'sp4_h_r_32')
// (8, 5, 'local_g1_7')
// (8, 5, 'lutff_1/in_3')
// (8, 5, 'sp12_h_r_23')
// (8, 5, 'sp4_h_r_45')
// (8, 6, 'local_g3_5')
// (8, 6, 'lutff_0/in_0')
// (8, 6, 'sp4_r_v_b_45')
// (8, 7, 'sp4_r_v_b_32')
// (8, 8, 'sp4_r_v_b_21')
// (8, 9, 'sp4_r_v_b_8')
// (9, 5, 'sp12_h_l_23')
// (9, 5, 'sp4_h_l_45')
// (9, 5, 'sp4_v_t_45')
// (9, 6, 'sp4_v_b_45')
// (9, 7, 'sp4_v_b_32')
// (9, 8, 'sp4_v_b_21')
// (9, 9, 'sp4_v_b_8')

wire n16;
// (0, 6, 'span12_horz_12')
// (1, 6, 'sp12_h_r_15')
// (2, 6, 'local_g1_0')
// (2, 6, 'lutff_3/in_2')
// (2, 6, 'sp12_h_r_16')
// (3, 5, 'neigh_op_tnr_6')
// (3, 6, 'neigh_op_rgt_6')
// (3, 6, 'sp12_h_r_19')
// (3, 7, 'neigh_op_bnr_6')
// (4, 5, 'neigh_op_top_6')
// (4, 6, 'local_g0_6')
// (4, 6, 'lutff_2/in_2')
// (4, 6, 'lutff_6/out')
// (4, 6, 'sp12_h_r_20')
// (4, 7, 'neigh_op_bot_6')
// (5, 5, 'neigh_op_tnl_6')
// (5, 6, 'neigh_op_lft_6')
// (5, 6, 'sp12_h_r_23')
// (5, 7, 'neigh_op_bnl_6')
// (6, 6, 'sp12_h_l_23')

reg n17 = 0;
// (0, 6, 'span12_horz_14')
// (1, 5, 'sp4_h_r_4')
// (1, 6, 'sp12_h_r_17')
// (1, 7, 'sp4_h_r_7')
// (2, 5, 'local_g0_1')
// (2, 5, 'lutff_0/in_1')
// (2, 5, 'sp4_h_r_17')
// (2, 6, 'local_g0_2')
// (2, 6, 'lutff_1/in_1')
// (2, 6, 'lutff_7/in_3')
// (2, 6, 'sp12_h_r_18')
// (2, 7, 'local_g0_2')
// (2, 7, 'lutff_0/in_2')
// (2, 7, 'lutff_4/in_2')
// (2, 7, 'lutff_7/in_3')
// (2, 7, 'sp4_h_r_18')
// (3, 5, 'neigh_op_tnr_7')
// (3, 5, 'sp4_h_r_28')
// (3, 6, 'neigh_op_rgt_7')
// (3, 6, 'sp12_h_r_21')
// (3, 7, 'neigh_op_bnr_7')
// (3, 7, 'sp4_h_r_31')
// (4, 4, 'sp4_r_v_b_39')
// (4, 5, 'neigh_op_top_7')
// (4, 5, 'sp4_h_r_41')
// (4, 5, 'sp4_r_v_b_26')
// (4, 6, 'local_g1_7')
// (4, 6, 'lutff_7/in_3')
// (4, 6, 'lutff_7/out')
// (4, 6, 'sp12_h_r_22')
// (4, 6, 'sp4_r_v_b_15')
// (4, 6, 'sp4_r_v_b_47')
// (4, 7, 'neigh_op_bot_7')
// (4, 7, 'sp4_h_r_42')
// (4, 7, 'sp4_r_v_b_2')
// (4, 7, 'sp4_r_v_b_34')
// (4, 8, 'sp4_r_v_b_23')
// (4, 9, 'sp4_r_v_b_10')
// (5, 3, 'sp4_v_t_39')
// (5, 4, 'sp4_v_b_39')
// (5, 5, 'neigh_op_tnl_7')
// (5, 5, 'sp4_h_l_41')
// (5, 5, 'sp4_v_b_26')
// (5, 5, 'sp4_v_t_47')
// (5, 6, 'neigh_op_lft_7')
// (5, 6, 'sp12_h_l_22')
// (5, 6, 'sp4_v_b_15')
// (5, 6, 'sp4_v_b_47')
// (5, 7, 'neigh_op_bnl_7')
// (5, 7, 'sp4_h_l_42')
// (5, 7, 'sp4_v_b_2')
// (5, 7, 'sp4_v_b_34')
// (5, 8, 'sp4_v_b_23')
// (5, 9, 'sp4_v_b_10')

wire n18;
// (0, 6, 'span12_horz_9')
// (1, 6, 'sp12_h_r_10')
// (2, 6, 'local_g1_5')
// (2, 6, 'lutff_3/in_1')
// (2, 6, 'sp12_h_r_13')
// (3, 6, 'sp12_h_r_14')
// (4, 5, 'neigh_op_tnr_5')
// (4, 6, 'local_g3_5')
// (4, 6, 'lutff_3/in_3')
// (4, 6, 'neigh_op_rgt_5')
// (4, 6, 'sp12_h_r_17')
// (4, 7, 'neigh_op_bnr_5')
// (5, 5, 'neigh_op_top_5')
// (5, 6, 'lutff_5/out')
// (5, 6, 'sp12_h_r_18')
// (5, 7, 'neigh_op_bot_5')
// (6, 5, 'neigh_op_tnl_5')
// (6, 6, 'neigh_op_lft_5')
// (6, 6, 'sp12_h_r_21')
// (6, 7, 'neigh_op_bnl_5')
// (7, 6, 'sp12_h_r_22')
// (8, 6, 'sp12_h_l_22')

reg d_vld = 0;
// (0, 7, 'logic_op_tnr_6')
// (0, 8, 'logic_op_rgt_6')
// (0, 9, 'logic_op_bnr_6')
// (0, 14, 'io_0/D_OUT_0')
// (0, 14, 'io_0/PAD')
// (0, 14, 'local_g1_7')
// (0, 14, 'span12_horz_23')
// (1, 2, 'sp12_v_t_23')
// (1, 3, 'sp12_v_b_23')
// (1, 4, 'sp12_v_b_20')
// (1, 5, 'sp12_v_b_19')
// (1, 6, 'sp12_v_b_16')
// (1, 7, 'neigh_op_top_6')
// (1, 7, 'sp12_v_b_15')
// (1, 8, 'lutff_6/out')
// (1, 8, 'sp12_v_b_12')
// (1, 9, 'neigh_op_bot_6')
// (1, 9, 'sp12_v_b_11')
// (1, 10, 'sp12_v_b_8')
// (1, 11, 'sp12_v_b_7')
// (1, 12, 'sp12_v_b_4')
// (1, 13, 'sp12_v_b_3')
// (1, 14, 'sp12_h_l_23')
// (1, 14, 'sp12_v_b_0')
// (2, 7, 'neigh_op_tnl_6')
// (2, 8, 'neigh_op_lft_6')
// (2, 9, 'neigh_op_bnl_6')

wire n20;
// (0, 7, 'span12_horz_2')
// (1, 7, 'sp12_h_r_5')
// (2, 7, 'sp12_h_r_6')
// (3, 6, 'neigh_op_tnr_1')
// (3, 7, 'neigh_op_rgt_1')
// (3, 7, 'sp12_h_r_9')
// (3, 8, 'neigh_op_bnr_1')
// (4, 5, 'sp4_r_v_b_43')
// (4, 6, 'neigh_op_top_1')
// (4, 6, 'sp4_r_v_b_30')
// (4, 7, 'lutff_1/out')
// (4, 7, 'sp12_h_r_10')
// (4, 7, 'sp4_r_v_b_19')
// (4, 8, 'neigh_op_bot_1')
// (4, 8, 'sp4_r_v_b_6')
// (5, 4, 'sp4_v_t_43')
// (5, 5, 'sp4_v_b_43')
// (5, 6, 'neigh_op_tnl_1')
// (5, 6, 'sp4_v_b_30')
// (5, 7, 'neigh_op_lft_1')
// (5, 7, 'sp12_h_r_13')
// (5, 7, 'sp4_v_b_19')
// (5, 8, 'local_g1_0')
// (5, 8, 'lutff_5/in_2')
// (5, 8, 'neigh_op_bnl_1')
// (5, 8, 'sp4_h_r_0')
// (5, 8, 'sp4_v_b_6')
// (6, 7, 'local_g1_6')
// (6, 7, 'lutff_5/in_2')
// (6, 7, 'sp12_h_r_14')
// (6, 8, 'sp4_h_r_13')
// (7, 7, 'sp12_h_r_17')
// (7, 8, 'sp4_h_r_24')
// (8, 7, 'sp12_h_r_18')
// (8, 8, 'sp4_h_r_37')
// (9, 7, 'sp12_h_r_21')
// (9, 8, 'sp4_h_l_37')
// (10, 7, 'sp12_h_r_22')
// (11, 7, 'sp12_h_l_22')

reg n21 = 0;
// (0, 7, 'span4_horz_4')
// (1, 6, 'neigh_op_tnr_6')
// (1, 7, 'neigh_op_rgt_6')
// (1, 7, 'sp4_h_r_17')
// (1, 7, 'sp4_r_v_b_44')
// (1, 8, 'neigh_op_bnr_6')
// (1, 8, 'sp4_r_v_b_33')
// (1, 9, 'sp4_r_v_b_20')
// (1, 10, 'sp4_r_v_b_9')
// (2, 1, 'sp12_v_t_23')
// (2, 2, 'sp12_v_b_23')
// (2, 3, 'sp12_v_b_20')
// (2, 4, 'sp12_v_b_19')
// (2, 5, 'sp12_v_b_16')
// (2, 6, 'neigh_op_top_6')
// (2, 6, 'sp12_v_b_15')
// (2, 6, 'sp4_v_t_44')
// (2, 7, 'lutff_6/out')
// (2, 7, 'sp12_v_b_12')
// (2, 7, 'sp4_h_r_28')
// (2, 7, 'sp4_v_b_44')
// (2, 8, 'neigh_op_bot_6')
// (2, 8, 'sp12_v_b_11')
// (2, 8, 'sp4_v_b_33')
// (2, 9, 'local_g2_0')
// (2, 9, 'local_g3_0')
// (2, 9, 'lutff_2/in_3')
// (2, 9, 'lutff_4/in_3')
// (2, 9, 'lutff_7/in_3')
// (2, 9, 'sp12_v_b_8')
// (2, 9, 'sp4_v_b_20')
// (2, 10, 'sp12_v_b_7')
// (2, 10, 'sp4_h_r_9')
// (2, 10, 'sp4_v_b_9')
// (2, 11, 'sp12_v_b_4')
// (2, 12, 'sp12_v_b_3')
// (2, 13, 'sp12_v_b_0')
// (3, 6, 'neigh_op_tnl_6')
// (3, 7, 'neigh_op_lft_6')
// (3, 7, 'sp4_h_r_41')
// (3, 8, 'neigh_op_bnl_6')
// (3, 8, 'sp4_r_v_b_41')
// (3, 8, 'sp4_r_v_b_44')
// (3, 9, 'sp4_r_v_b_28')
// (3, 9, 'sp4_r_v_b_33')
// (3, 10, 'sp4_h_r_20')
// (3, 10, 'sp4_r_v_b_17')
// (3, 10, 'sp4_r_v_b_20')
// (3, 11, 'sp4_r_v_b_4')
// (3, 11, 'sp4_r_v_b_9')
// (4, 7, 'sp4_h_l_41')
// (4, 7, 'sp4_h_r_3')
// (4, 7, 'sp4_v_t_41')
// (4, 7, 'sp4_v_t_44')
// (4, 8, 'local_g2_4')
// (4, 8, 'lutff_1/in_3')
// (4, 8, 'sp4_v_b_41')
// (4, 8, 'sp4_v_b_44')
// (4, 9, 'sp4_v_b_28')
// (4, 9, 'sp4_v_b_33')
// (4, 10, 'local_g1_1')
// (4, 10, 'local_g2_1')
// (4, 10, 'lutff_1/in_3')
// (4, 10, 'lutff_6/in_3')
// (4, 10, 'lutff_7/in_3')
// (4, 10, 'sp4_h_r_33')
// (4, 10, 'sp4_v_b_17')
// (4, 10, 'sp4_v_b_20')
// (4, 11, 'local_g1_1')
// (4, 11, 'local_g1_4')
// (4, 11, 'lutff_1/in_3')
// (4, 11, 'lutff_2/in_3')
// (4, 11, 'lutff_4/in_3')
// (4, 11, 'sp4_h_r_9')
// (4, 11, 'sp4_v_b_4')
// (4, 11, 'sp4_v_b_9')
// (5, 7, 'sp4_h_r_14')
// (5, 7, 'sp4_r_v_b_38')
// (5, 7, 'sp4_r_v_b_39')
// (5, 8, 'sp4_r_v_b_26')
// (5, 8, 'sp4_r_v_b_27')
// (5, 9, 'sp4_r_v_b_14')
// (5, 9, 'sp4_r_v_b_15')
// (5, 10, 'sp4_h_r_44')
// (5, 10, 'sp4_r_v_b_2')
// (5, 10, 'sp4_r_v_b_3')
// (5, 11, 'sp4_h_r_20')
// (6, 6, 'sp4_v_t_38')
// (6, 6, 'sp4_v_t_39')
// (6, 7, 'sp4_h_r_27')
// (6, 7, 'sp4_v_b_38')
// (6, 7, 'sp4_v_b_39')
// (6, 8, 'sp4_v_b_26')
// (6, 8, 'sp4_v_b_27')
// (6, 9, 'local_g0_6')
// (6, 9, 'local_g1_6')
// (6, 9, 'lutff_1/in_3')
// (6, 9, 'lutff_3/in_3')
// (6, 9, 'lutff_6/in_3')
// (6, 9, 'sp4_v_b_14')
// (6, 9, 'sp4_v_b_15')
// (6, 10, 'local_g0_2')
// (6, 10, 'local_g0_3')
// (6, 10, 'lutff_0/in_3')
// (6, 10, 'lutff_3/in_3')
// (6, 10, 'lutff_5/in_3')
// (6, 10, 'sp4_h_l_44')
// (6, 10, 'sp4_h_r_9')
// (6, 10, 'sp4_v_b_2')
// (6, 10, 'sp4_v_b_3')
// (6, 11, 'local_g2_1')
// (6, 11, 'local_g3_1')
// (6, 11, 'lutff_0/in_3')
// (6, 11, 'lutff_3/in_3')
// (6, 11, 'lutff_5/in_3')
// (6, 11, 'sp4_h_r_33')
// (7, 7, 'sp4_h_r_38')
// (7, 8, 'local_g3_4')
// (7, 8, 'local_g3_5')
// (7, 8, 'lutff_0/in_3')
// (7, 8, 'lutff_6/in_3')
// (7, 8, 'lutff_7/in_3')
// (7, 8, 'sp4_r_v_b_44')
// (7, 8, 'sp4_r_v_b_45')
// (7, 9, 'sp4_r_v_b_32')
// (7, 9, 'sp4_r_v_b_33')
// (7, 10, 'local_g0_4')
// (7, 10, 'local_g3_4')
// (7, 10, 'lutff_0/in_3')
// (7, 10, 'lutff_4/in_3')
// (7, 10, 'lutff_7/in_3')
// (7, 10, 'sp4_h_r_20')
// (7, 10, 'sp4_r_v_b_20')
// (7, 10, 'sp4_r_v_b_21')
// (7, 11, 'sp4_h_r_44')
// (7, 11, 'sp4_r_v_b_8')
// (7, 11, 'sp4_r_v_b_9')
// (8, 7, 'sp4_h_l_38')
// (8, 7, 'sp4_v_t_44')
// (8, 7, 'sp4_v_t_45')
// (8, 8, 'sp4_v_b_44')
// (8, 8, 'sp4_v_b_45')
// (8, 9, 'sp4_v_b_32')
// (8, 9, 'sp4_v_b_33')
// (8, 10, 'sp4_h_r_33')
// (8, 10, 'sp4_v_b_20')
// (8, 10, 'sp4_v_b_21')
// (8, 11, 'sp4_h_l_44')
// (8, 11, 'sp4_v_b_8')
// (8, 11, 'sp4_v_b_9')
// (9, 10, 'sp4_h_r_44')
// (10, 10, 'sp4_h_l_44')

wire n22;
// (0, 8, 'span12_horz_12')
// (1, 8, 'sp12_h_r_15')
// (2, 8, 'local_g1_0')
// (2, 8, 'lutff_2/in_3')
// (2, 8, 'sp12_h_r_0')
// (2, 8, 'sp12_h_r_16')
// (3, 7, 'neigh_op_tnr_6')
// (3, 8, 'neigh_op_rgt_6')
// (3, 8, 'sp12_h_r_19')
// (3, 8, 'sp12_h_r_3')
// (3, 9, 'neigh_op_bnr_6')
// (4, 7, 'neigh_op_top_6')
// (4, 8, 'lutff_6/out')
// (4, 8, 'sp12_h_r_20')
// (4, 8, 'sp12_h_r_4')
// (4, 9, 'neigh_op_bot_6')
// (5, 7, 'neigh_op_tnl_6')
// (5, 8, 'neigh_op_lft_6')
// (5, 8, 'sp12_h_r_23')
// (5, 8, 'sp12_h_r_7')
// (5, 9, 'neigh_op_bnl_6')
// (6, 8, 'sp12_h_l_23')
// (6, 8, 'sp12_h_r_8')
// (7, 8, 'local_g0_3')
// (7, 8, 'local_g1_3')
// (7, 8, 'lutff_1/in_3')
// (7, 8, 'lutff_4/in_3')
// (7, 8, 'sp12_h_r_11')
// (8, 8, 'sp12_h_r_12')
// (9, 8, 'sp12_h_r_15')
// (10, 8, 'sp12_h_r_16')
// (11, 8, 'sp12_h_r_19')
// (12, 8, 'sp12_h_r_20')
// (13, 8, 'span12_horz_20')

reg n23 = 0;
// (0, 8, 'span12_horz_2')
// (1, 8, 'sp12_h_r_5')
// (2, 8, 'sp12_h_r_6')
// (3, 8, 'sp12_h_r_9')
// (4, 8, 'sp12_h_r_10')
// (5, 7, 'neigh_op_tnr_3')
// (5, 8, 'local_g2_3')
// (5, 8, 'lutff_7/in_0')
// (5, 8, 'neigh_op_rgt_3')
// (5, 8, 'sp12_h_r_13')
// (5, 9, 'neigh_op_bnr_3')
// (6, 7, 'neigh_op_top_3')
// (6, 8, 'lutff_3/out')
// (6, 8, 'sp12_h_r_14')
// (6, 9, 'neigh_op_bot_3')
// (7, 7, 'neigh_op_tnl_3')
// (7, 8, 'local_g0_1')
// (7, 8, 'lutff_4/in_1')
// (7, 8, 'neigh_op_lft_3')
// (7, 8, 'sp12_h_r_17')
// (7, 9, 'neigh_op_bnl_3')
// (8, 8, 'sp12_h_r_18')
// (9, 8, 'sp12_h_r_21')
// (10, 8, 'sp12_h_r_22')
// (11, 8, 'sp12_h_l_22')

reg n24 = 0;
// (0, 8, 'span12_horz_6')
// (1, 8, 'sp12_h_r_9')
// (2, 8, 'sp12_h_r_10')
// (3, 8, 'sp12_h_r_13')
// (4, 8, 'sp12_h_r_14')
// (5, 7, 'neigh_op_tnr_5')
// (5, 8, 'neigh_op_rgt_5')
// (5, 8, 'sp12_h_r_17')
// (5, 9, 'neigh_op_bnr_5')
// (6, 7, 'neigh_op_top_5')
// (6, 8, 'local_g0_2')
// (6, 8, 'lutff_4/in_0')
// (6, 8, 'lutff_5/out')
// (6, 8, 'sp12_h_r_18')
// (6, 9, 'neigh_op_bot_5')
// (7, 7, 'neigh_op_tnl_5')
// (7, 8, 'neigh_op_lft_5')
// (7, 8, 'sp12_h_r_21')
// (7, 9, 'neigh_op_bnl_5')
// (8, 8, 'sp12_h_r_22')
// (9, 8, 'sp12_h_l_22')

wire n25;
// (0, 8, 'span12_horz_8')
// (1, 8, 'sp12_h_r_11')
// (2, 8, 'sp12_h_r_12')
// (2, 8, 'sp4_h_r_0')
// (3, 5, 'sp4_r_v_b_45')
// (3, 6, 'sp4_r_v_b_32')
// (3, 7, 'neigh_op_tnr_4')
// (3, 7, 'sp4_r_v_b_21')
// (3, 8, 'neigh_op_rgt_4')
// (3, 8, 'sp12_h_r_15')
// (3, 8, 'sp4_h_r_13')
// (3, 8, 'sp4_r_v_b_8')
// (3, 9, 'neigh_op_bnr_4')
// (4, 4, 'sp4_v_t_45')
// (4, 5, 'local_g3_5')
// (4, 5, 'lutff_5/in_3')
// (4, 5, 'sp4_v_b_45')
// (4, 6, 'sp4_v_b_32')
// (4, 7, 'neigh_op_top_4')
// (4, 7, 'sp4_v_b_21')
// (4, 8, 'lutff_4/out')
// (4, 8, 'sp12_h_r_16')
// (4, 8, 'sp4_h_r_2')
// (4, 8, 'sp4_h_r_24')
// (4, 8, 'sp4_v_b_8')
// (4, 9, 'local_g1_4')
// (4, 9, 'lutff_5/in_2')
// (4, 9, 'neigh_op_bot_4')
// (5, 7, 'neigh_op_tnl_4')
// (5, 8, 'neigh_op_lft_4')
// (5, 8, 'sp12_h_r_19')
// (5, 8, 'sp4_h_r_15')
// (5, 8, 'sp4_h_r_37')
// (5, 9, 'neigh_op_bnl_4')
// (5, 9, 'sp4_r_v_b_37')
// (5, 10, 'sp4_r_v_b_24')
// (5, 11, 'sp4_r_v_b_13')
// (5, 12, 'sp4_r_v_b_0')
// (6, 8, 'local_g1_4')
// (6, 8, 'lutff_0/in_3')
// (6, 8, 'sp12_h_r_20')
// (6, 8, 'sp4_h_l_37')
// (6, 8, 'sp4_h_r_26')
// (6, 8, 'sp4_v_t_37')
// (6, 9, 'local_g2_5')
// (6, 9, 'local_g3_5')
// (6, 9, 'lutff_4/in_3')
// (6, 9, 'lutff_7/in_3')
// (6, 9, 'sp4_v_b_37')
// (6, 10, 'local_g2_0')
// (6, 10, 'lutff_7/in_3')
// (6, 10, 'sp4_v_b_24')
// (6, 11, 'sp4_v_b_13')
// (6, 12, 'sp4_v_b_0')
// (7, 8, 'local_g0_7')
// (7, 8, 'lutff_1/in_2')
// (7, 8, 'sp12_h_r_23')
// (7, 8, 'sp4_h_r_39')
// (7, 9, 'sp4_r_v_b_39')
// (7, 10, 'local_g0_2')
// (7, 10, 'lutff_1/in_3')
// (7, 10, 'sp4_r_v_b_26')
// (7, 11, 'sp4_r_v_b_15')
// (7, 12, 'sp4_r_v_b_2')
// (8, 8, 'sp12_h_l_23')
// (8, 8, 'sp4_h_l_39')
// (8, 8, 'sp4_v_t_39')
// (8, 9, 'sp4_v_b_39')
// (8, 10, 'sp4_v_b_26')
// (8, 11, 'sp4_v_b_15')
// (8, 12, 'sp4_v_b_2')

reg n26 = 0;
// (0, 9, 'span12_horz_1')
// (1, 9, 'sp12_h_r_2')
// (2, 9, 'sp12_h_r_5')
// (3, 9, 'sp12_h_r_6')
// (4, 9, 'sp12_h_r_9')
// (5, 9, 'sp12_h_r_10')
// (6, 9, 'sp12_h_r_13')
// (7, 9, 'sp12_h_r_14')
// (8, 9, 'local_g1_1')
// (8, 9, 'lutff_1/in_1')
// (8, 9, 'lutff_3/in_1')
// (8, 9, 'sp12_h_r_17')
// (9, 9, 'sp12_h_r_18')
// (10, 8, 'neigh_op_tnr_7')
// (10, 9, 'neigh_op_rgt_7')
// (10, 9, 'sp12_h_r_21')
// (10, 10, 'neigh_op_bnr_7')
// (11, 8, 'neigh_op_top_7')
// (11, 9, 'lutff_7/out')
// (11, 9, 'sp12_h_r_22')
// (11, 10, 'neigh_op_bot_7')
// (12, 8, 'neigh_op_tnl_7')
// (12, 9, 'neigh_op_lft_7')
// (12, 9, 'sp12_h_l_22')
// (12, 10, 'neigh_op_bnl_7')

reg n27 = 0;
// (0, 10, 'span12_horz_3')
// (1, 10, 'sp12_h_r_4')
// (2, 10, 'sp12_h_r_7')
// (3, 10, 'sp12_h_r_8')
// (4, 9, 'neigh_op_tnr_2')
// (4, 10, 'neigh_op_rgt_2')
// (4, 10, 'sp12_h_r_11')
// (4, 11, 'neigh_op_bnr_2')
// (5, 9, 'neigh_op_top_2')
// (5, 10, 'lutff_2/out')
// (5, 10, 'sp12_h_r_12')
// (5, 11, 'neigh_op_bot_2')
// (6, 9, 'neigh_op_tnl_2')
// (6, 10, 'neigh_op_lft_2')
// (6, 10, 'sp12_h_r_15')
// (6, 11, 'neigh_op_bnl_2')
// (7, 10, 'local_g0_0')
// (7, 10, 'lutff_7/in_1')
// (7, 10, 'sp12_h_r_16')
// (8, 10, 'sp12_h_r_19')
// (9, 10, 'sp12_h_r_20')
// (10, 10, 'sp12_h_r_23')
// (11, 10, 'sp12_h_l_23')

reg n28 = 0;
// (0, 10, 'span12_horz_4')
// (1, 10, 'sp12_h_r_7')
// (2, 10, 'sp12_h_r_8')
// (3, 9, 'neigh_op_tnr_2')
// (3, 10, 'neigh_op_rgt_2')
// (3, 10, 'sp12_h_r_11')
// (3, 11, 'neigh_op_bnr_2')
// (4, 9, 'neigh_op_top_2')
// (4, 10, 'local_g0_2')
// (4, 10, 'local_g1_4')
// (4, 10, 'lutff_2/out')
// (4, 10, 'lutff_3/in_1')
// (4, 10, 'lutff_7/in_2')
// (4, 10, 'sp12_h_r_12')
// (4, 11, 'neigh_op_bot_2')
// (5, 9, 'neigh_op_tnl_2')
// (5, 10, 'neigh_op_lft_2')
// (5, 10, 'sp12_h_r_15')
// (5, 11, 'neigh_op_bnl_2')
// (6, 10, 'sp12_h_r_16')
// (7, 10, 'sp12_h_r_19')
// (8, 10, 'sp12_h_r_20')
// (9, 10, 'sp12_h_r_23')
// (10, 10, 'sp12_h_l_23')

reg n29 = 0;
// (0, 10, 'span4_horz_2')
// (1, 10, 'sp4_h_r_15')
// (2, 10, 'local_g2_2')
// (2, 10, 'lutff_2/in_0')
// (2, 10, 'sp4_h_r_26')
// (3, 7, 'sp4_r_v_b_44')
// (3, 8, 'neigh_op_tnr_2')
// (3, 8, 'sp4_r_v_b_33')
// (3, 9, 'neigh_op_rgt_2')
// (3, 9, 'sp4_r_v_b_20')
// (3, 10, 'neigh_op_bnr_2')
// (3, 10, 'sp4_h_r_39')
// (3, 10, 'sp4_r_v_b_9')
// (4, 6, 'sp4_v_t_44')
// (4, 7, 'sp4_v_b_44')
// (4, 8, 'neigh_op_top_2')
// (4, 8, 'sp4_v_b_33')
// (4, 9, 'lutff_2/out')
// (4, 9, 'sp4_v_b_20')
// (4, 10, 'local_g0_1')
// (4, 10, 'lutff_2/in_1')
// (4, 10, 'neigh_op_bot_2')
// (4, 10, 'sp4_h_l_39')
// (4, 10, 'sp4_v_b_9')
// (5, 8, 'neigh_op_tnl_2')
// (5, 9, 'neigh_op_lft_2')
// (5, 10, 'neigh_op_bnl_2')

reg n30 = 0;
// (0, 11, 'span12_horz_8')
// (1, 10, 'neigh_op_tnr_2')
// (1, 11, 'neigh_op_rgt_2')
// (1, 11, 'sp12_h_r_11')
// (1, 12, 'neigh_op_bnr_2')
// (2, 9, 'sp12_h_r_0')
// (2, 9, 'sp12_v_t_23')
// (2, 10, 'neigh_op_top_2')
// (2, 10, 'sp12_v_b_23')
// (2, 11, 'lutff_2/out')
// (2, 11, 'sp12_h_r_12')
// (2, 11, 'sp12_v_b_20')
// (2, 12, 'neigh_op_bot_2')
// (2, 12, 'sp12_v_b_19')
// (2, 13, 'sp12_v_b_16')
// (2, 14, 'sp12_v_b_15')
// (2, 15, 'sp12_v_b_12')
// (2, 16, 'sp12_v_b_11')
// (2, 17, 'span12_vert_8')
// (3, 9, 'sp12_h_r_3')
// (3, 10, 'neigh_op_tnl_2')
// (3, 11, 'neigh_op_lft_2')
// (3, 11, 'sp12_h_r_15')
// (3, 12, 'neigh_op_bnl_2')
// (4, 9, 'sp12_h_r_4')
// (4, 11, 'sp12_h_r_16')
// (5, 9, 'sp12_h_r_7')
// (5, 11, 'local_g1_3')
// (5, 11, 'lutff_6/in_0')
// (5, 11, 'sp12_h_r_19')
// (6, 9, 'sp12_h_r_8')
// (6, 11, 'sp12_h_r_20')
// (7, 9, 'local_g1_3')
// (7, 9, 'lutff_2/in_0')
// (7, 9, 'lutff_6/in_0')
// (7, 9, 'sp12_h_r_11')
// (7, 11, 'local_g0_7')
// (7, 11, 'lutff_7/in_0')
// (7, 11, 'sp12_h_r_23')
// (8, 9, 'sp12_h_r_12')
// (8, 11, 'sp12_h_l_23')
// (9, 9, 'sp12_h_r_15')
// (10, 9, 'sp12_h_r_16')
// (11, 9, 'sp12_h_r_19')
// (12, 9, 'sp12_h_r_20')
// (13, 9, 'span12_horz_20')

reg n31 = 0;
// (0, 12, 'span12_horz_2')
// (1, 11, 'neigh_op_tnr_7')
// (1, 12, 'neigh_op_rgt_7')
// (1, 12, 'sp12_h_r_5')
// (1, 13, 'neigh_op_bnr_7')
// (2, 11, 'neigh_op_top_7')
// (2, 12, 'lutff_7/out')
// (2, 12, 'sp12_h_r_6')
// (2, 13, 'neigh_op_bot_7')
// (3, 11, 'neigh_op_tnl_7')
// (3, 12, 'neigh_op_lft_7')
// (3, 12, 'sp12_h_r_9')
// (3, 13, 'neigh_op_bnl_7')
// (4, 12, 'local_g1_2')
// (4, 12, 'lutff_1/in_0')
// (4, 12, 'sp12_h_r_10')
// (5, 12, 'sp12_h_r_13')
// (6, 12, 'sp12_h_r_14')
// (7, 12, 'sp12_h_r_17')
// (8, 12, 'sp12_h_r_18')
// (9, 12, 'sp12_h_r_21')
// (10, 12, 'sp12_h_r_22')
// (11, 12, 'sp12_h_l_22')

reg n32 = 0;
// (0, 13, 'span12_horz_0')
// (1, 13, 'sp12_h_r_3')
// (2, 13, 'sp12_h_r_4')
// (3, 13, 'sp12_h_r_7')
// (4, 13, 'sp12_h_r_8')
// (5, 13, 'sp12_h_r_11')
// (6, 13, 'sp12_h_r_12')
// (7, 12, 'neigh_op_tnr_4')
// (7, 13, 'neigh_op_rgt_4')
// (7, 13, 'sp12_h_r_15')
// (7, 14, 'neigh_op_bnr_4')
// (8, 12, 'neigh_op_top_4')
// (8, 13, 'lutff_4/out')
// (8, 13, 'sp12_h_r_16')
// (8, 14, 'neigh_op_bot_4')
// (9, 12, 'neigh_op_tnl_4')
// (9, 13, 'neigh_op_lft_4')
// (9, 13, 'sp12_h_r_19')
// (9, 14, 'neigh_op_bnl_4')
// (10, 13, 'sp12_h_r_20')
// (11, 13, 'local_g0_7')
// (11, 13, 'lutff_5/in_0')
// (11, 13, 'sp12_h_r_23')
// (12, 13, 'sp12_h_l_23')

reg n33 = 0;
// (0, 13, 'span12_horz_10')
// (1, 13, 'sp12_h_r_13')
// (2, 13, 'sp12_h_r_14')
// (3, 13, 'sp12_h_r_17')
// (4, 13, 'sp12_h_r_18')
// (5, 13, 'sp12_h_r_21')
// (6, 13, 'local_g1_6')
// (6, 13, 'lutff_7/in_0')
// (6, 13, 'sp12_h_r_22')
// (7, 12, 'neigh_op_tnr_5')
// (7, 13, 'neigh_op_rgt_5')
// (7, 13, 'sp12_h_l_22')
// (7, 13, 'sp12_h_r_1')
// (7, 14, 'neigh_op_bnr_5')
// (8, 12, 'neigh_op_top_5')
// (8, 13, 'lutff_5/out')
// (8, 13, 'sp12_h_r_2')
// (8, 14, 'neigh_op_bot_5')
// (9, 12, 'neigh_op_tnl_5')
// (9, 13, 'neigh_op_lft_5')
// (9, 13, 'sp12_h_r_5')
// (9, 14, 'neigh_op_bnl_5')
// (10, 13, 'sp12_h_r_6')
// (11, 13, 'sp12_h_r_9')
// (12, 13, 'sp12_h_r_10')
// (13, 13, 'span12_horz_10')

reg n34 = 0;
// (0, 13, 'span12_horz_14')
// (1, 13, 'sp12_h_r_17')
// (2, 13, 'local_g0_2')
// (2, 13, 'lutff_0/in_0')
// (2, 13, 'sp12_h_r_18')
// (3, 12, 'neigh_op_tnr_7')
// (3, 13, 'neigh_op_rgt_7')
// (3, 13, 'sp12_h_r_21')
// (3, 14, 'neigh_op_bnr_7')
// (4, 12, 'neigh_op_top_7')
// (4, 13, 'local_g0_7')
// (4, 13, 'lutff_5/in_0')
// (4, 13, 'lutff_7/out')
// (4, 13, 'sp12_h_r_22')
// (4, 14, 'neigh_op_bot_7')
// (5, 12, 'local_g2_7')
// (5, 12, 'local_g3_7')
// (5, 12, 'lutff_1/in_0')
// (5, 12, 'lutff_6/in_0')
// (5, 12, 'neigh_op_tnl_7')
// (5, 13, 'neigh_op_lft_7')
// (5, 13, 'sp12_h_l_22')
// (5, 14, 'neigh_op_bnl_7')

reg n35 = 0;
// (0, 13, 'span12_horz_2')
// (1, 13, 'sp12_h_r_5')
// (2, 13, 'local_g1_6')
// (2, 13, 'lutff_3/in_0')
// (2, 13, 'sp12_h_r_6')
// (3, 13, 'sp12_h_r_9')
// (4, 13, 'sp12_h_r_10')
// (5, 12, 'neigh_op_tnr_3')
// (5, 13, 'neigh_op_rgt_3')
// (5, 13, 'sp12_h_r_13')
// (5, 14, 'neigh_op_bnr_3')
// (6, 12, 'neigh_op_top_3')
// (6, 13, 'lutff_3/out')
// (6, 13, 'sp12_h_r_14')
// (6, 14, 'neigh_op_bot_3')
// (7, 12, 'neigh_op_tnl_3')
// (7, 13, 'neigh_op_lft_3')
// (7, 13, 'sp12_h_r_17')
// (7, 14, 'neigh_op_bnl_3')
// (8, 13, 'sp12_h_r_18')
// (9, 13, 'sp12_h_r_21')
// (10, 13, 'sp12_h_r_22')
// (11, 13, 'sp12_h_l_22')

reg n36 = 0;
// (0, 13, 'span12_horz_5')
// (1, 13, 'sp12_h_r_6')
// (2, 13, 'sp12_h_r_9')
// (3, 13, 'sp12_h_r_10')
// (4, 12, 'neigh_op_tnr_3')
// (4, 13, 'neigh_op_rgt_3')
// (4, 13, 'sp12_h_r_13')
// (4, 14, 'neigh_op_bnr_3')
// (5, 12, 'neigh_op_top_3')
// (5, 13, 'local_g0_6')
// (5, 13, 'lutff_2/in_0')
// (5, 13, 'lutff_3/out')
// (5, 13, 'sp12_h_r_14')
// (5, 14, 'neigh_op_bot_3')
// (6, 12, 'neigh_op_tnl_3')
// (6, 13, 'neigh_op_lft_3')
// (6, 13, 'sp12_h_r_17')
// (6, 14, 'neigh_op_bnl_3')
// (7, 13, 'sp12_h_r_18')
// (8, 13, 'sp12_h_r_21')
// (9, 13, 'sp12_h_r_22')
// (10, 13, 'sp12_h_l_22')

reg n37 = 0;
// (0, 13, 'span12_horz_8')
// (1, 13, 'sp12_h_r_11')
// (2, 13, 'local_g1_4')
// (2, 13, 'lutff_0/in_1')
// (2, 13, 'sp12_h_r_12')
// (3, 12, 'neigh_op_tnr_4')
// (3, 13, 'neigh_op_rgt_4')
// (3, 13, 'sp12_h_r_15')
// (3, 14, 'neigh_op_bnr_4')
// (4, 12, 'neigh_op_top_4')
// (4, 13, 'local_g1_4')
// (4, 13, 'lutff_0/in_1')
// (4, 13, 'lutff_4/out')
// (4, 13, 'sp12_h_r_16')
// (4, 14, 'neigh_op_bot_4')
// (5, 12, 'neigh_op_tnl_4')
// (5, 13, 'neigh_op_lft_4')
// (5, 13, 'sp12_h_r_19')
// (5, 14, 'neigh_op_bnl_4')
// (6, 13, 'sp12_h_r_20')
// (7, 13, 'sp12_h_r_23')
// (8, 13, 'sp12_h_l_23')

reg n38 = 0;
// (0, 13, 'span4_horz_0')
// (1, 12, 'neigh_op_tnr_4')
// (1, 13, 'neigh_op_rgt_4')
// (1, 13, 'sp4_h_r_13')
// (1, 14, 'neigh_op_bnr_4')
// (2, 12, 'neigh_op_top_4')
// (2, 13, 'lutff_4/out')
// (2, 13, 'sp4_h_r_24')
// (2, 14, 'neigh_op_bot_4')
// (3, 12, 'neigh_op_tnl_4')
// (3, 13, 'neigh_op_lft_4')
// (3, 13, 'sp4_h_r_37')
// (3, 14, 'neigh_op_bnl_4')
// (3, 14, 'sp4_r_v_b_40')
// (3, 15, 'sp4_r_v_b_29')
// (3, 16, 'sp4_r_v_b_16')
// (4, 13, 'sp4_h_l_37')
// (4, 13, 'sp4_v_t_40')
// (4, 14, 'local_g2_0')
// (4, 14, 'lutff_6/in_0')
// (4, 14, 'sp4_v_b_40')
// (4, 15, 'sp4_v_b_29')
// (4, 16, 'sp4_v_b_16')
// (4, 17, 'span4_vert_5')

wire rst;
// (0, 14, 'io_1/D_IN_0')
// (0, 14, 'io_1/PAD')
// (0, 14, 'span12_horz_20')
// (1, 2, 'sp4_h_r_1')
// (1, 7, 'sp4_r_v_b_41')
// (1, 8, 'local_g1_4')
// (1, 8, 'lutff_6/in_3')
// (1, 8, 'sp4_r_v_b_28')
// (1, 9, 'sp4_r_v_b_17')
// (1, 10, 'sp4_r_v_b_4')
// (1, 13, 'neigh_op_tnl_2')
// (1, 13, 'neigh_op_tnl_6')
// (1, 14, 'neigh_op_lft_2')
// (1, 14, 'neigh_op_lft_6')
// (1, 14, 'sp12_h_r_23')
// (1, 15, 'neigh_op_bnl_2')
// (1, 15, 'neigh_op_bnl_6')
// (2, 2, 'local_g1_0')
// (2, 2, 'lutff_4/in_3')
// (2, 2, 'lutff_6/in_1')
// (2, 2, 'sp12_h_r_0')
// (2, 2, 'sp12_v_t_23')
// (2, 2, 'sp4_h_r_12')
// (2, 3, 'sp12_v_b_23')
// (2, 4, 'sp12_v_b_20')
// (2, 5, 'sp12_v_b_19')
// (2, 6, 'local_g3_0')
// (2, 6, 'lutff_0/in_3')
// (2, 6, 'sp12_v_b_16')
// (2, 6, 'sp4_v_t_41')
// (2, 7, 'sp12_v_b_15')
// (2, 7, 'sp4_v_b_41')
// (2, 8, 'sp12_v_b_12')
// (2, 8, 'sp4_v_b_28')
// (2, 9, 'sp12_v_b_11')
// (2, 9, 'sp4_v_b_17')
// (2, 10, 'sp12_v_b_8')
// (2, 10, 'sp4_v_b_4')
// (2, 11, 'sp12_v_b_7')
// (2, 12, 'sp12_v_b_4')
// (2, 13, 'sp12_v_b_3')
// (2, 14, 'sp12_h_l_23')
// (2, 14, 'sp12_v_b_0')
// (3, 2, 'sp12_h_r_3')
// (3, 2, 'sp4_h_r_25')
// (4, 2, 'local_g2_4')
// (4, 2, 'local_g3_4')
// (4, 2, 'lutff_2/in_1')
// (4, 2, 'lutff_7/in_3')
// (4, 2, 'sp12_h_r_4')
// (4, 2, 'sp4_h_r_36')
// (4, 3, 'local_g2_4')
// (4, 3, 'lutff_global/s_r')
// (4, 3, 'sp4_r_v_b_36')
// (4, 4, 'sp4_r_v_b_25')
// (4, 5, 'sp4_r_v_b_12')
// (4, 6, 'sp4_r_v_b_1')
// (5, 2, 'local_g0_7')
// (5, 2, 'local_g1_7')
// (5, 2, 'lutff_3/in_3')
// (5, 2, 'lutff_5/in_3')
// (5, 2, 'lutff_6/in_3')
// (5, 2, 'lutff_7/in_3')
// (5, 2, 'sp12_h_r_7')
// (5, 2, 'sp4_h_l_36')
// (5, 2, 'sp4_v_t_36')
// (5, 3, 'sp4_v_b_36')
// (5, 4, 'sp4_v_b_25')
// (5, 5, 'sp4_v_b_12')
// (5, 6, 'sp4_v_b_1')
// (6, 2, 'sp12_h_r_8')
// (7, 2, 'sp12_h_r_11')
// (8, 2, 'sp12_h_r_12')
// (9, 2, 'sp12_h_r_15')
// (10, 2, 'sp12_h_r_16')
// (11, 2, 'sp12_h_r_19')
// (12, 2, 'sp12_h_r_20')
// (13, 2, 'span12_horz_20')

reg n40 = 0;
// (0, 14, 'span12_horz_6')
// (1, 14, 'sp12_h_r_9')
// (2, 14, 'local_g1_2')
// (2, 14, 'lutff_5/in_0')
// (2, 14, 'sp12_h_r_10')
// (3, 14, 'sp12_h_r_13')
// (4, 14, 'sp12_h_r_14')
// (5, 13, 'neigh_op_tnr_5')
// (5, 14, 'neigh_op_rgt_5')
// (5, 14, 'sp12_h_r_17')
// (5, 15, 'neigh_op_bnr_5')
// (6, 13, 'neigh_op_top_5')
// (6, 14, 'lutff_5/out')
// (6, 14, 'sp12_h_r_18')
// (6, 15, 'neigh_op_bot_5')
// (7, 13, 'neigh_op_tnl_5')
// (7, 14, 'neigh_op_lft_5')
// (7, 14, 'sp12_h_r_21')
// (7, 15, 'neigh_op_bnl_5')
// (8, 14, 'sp12_h_r_22')
// (9, 14, 'sp12_h_l_22')

reg n41 = 0;
// (1, 2, 'sp12_h_r_1')
// (2, 2, 'sp12_h_r_2')
// (3, 1, 'neigh_op_tnr_7')
// (3, 2, 'neigh_op_rgt_7')
// (3, 2, 'sp12_h_r_5')
// (3, 2, 'sp4_h_r_3')
// (3, 3, 'neigh_op_bnr_7')
// (4, 1, 'neigh_op_top_7')
// (4, 1, 'sp4_r_v_b_42')
// (4, 2, 'local_g1_7')
// (4, 2, 'lutff_1/in_3')
// (4, 2, 'lutff_7/in_1')
// (4, 2, 'lutff_7/out')
// (4, 2, 'sp12_h_r_6')
// (4, 2, 'sp4_h_r_14')
// (4, 2, 'sp4_r_v_b_31')
// (4, 3, 'neigh_op_bot_7')
// (4, 3, 'sp4_r_v_b_18')
// (4, 4, 'sp4_r_v_b_7')
// (5, 0, 'span4_vert_42')
// (5, 1, 'neigh_op_tnl_7')
// (5, 1, 'sp4_v_b_42')
// (5, 2, 'local_g0_1')
// (5, 2, 'lutff_6/in_1')
// (5, 2, 'neigh_op_lft_7')
// (5, 2, 'sp12_h_r_9')
// (5, 2, 'sp4_h_r_27')
// (5, 2, 'sp4_v_b_31')
// (5, 3, 'local_g2_7')
// (5, 3, 'lutff_3/in_2')
// (5, 3, 'neigh_op_bnl_7')
// (5, 3, 'sp4_v_b_18')
// (5, 4, 'local_g0_7')
// (5, 4, 'lutff_1/in_2')
// (5, 4, 'sp4_h_r_6')
// (5, 4, 'sp4_h_r_7')
// (5, 4, 'sp4_v_b_7')
// (6, 2, 'sp12_h_r_10')
// (6, 2, 'sp4_h_r_38')
// (6, 3, 'sp4_r_v_b_38')
// (6, 4, 'local_g1_3')
// (6, 4, 'lutff_3/in_3')
// (6, 4, 'sp4_h_r_18')
// (6, 4, 'sp4_h_r_19')
// (6, 4, 'sp4_r_v_b_27')
// (6, 5, 'sp4_r_v_b_14')
// (6, 6, 'sp4_r_v_b_3')
// (7, 2, 'sp12_h_r_13')
// (7, 2, 'sp4_h_l_38')
// (7, 2, 'sp4_h_r_8')
// (7, 2, 'sp4_v_t_38')
// (7, 3, 'sp4_v_b_38')
// (7, 4, 'local_g2_7')
// (7, 4, 'lutff_7/in_2')
// (7, 4, 'sp4_h_r_30')
// (7, 4, 'sp4_h_r_31')
// (7, 4, 'sp4_v_b_27')
// (7, 5, 'local_g0_6')
// (7, 5, 'lutff_4/in_2')
// (7, 5, 'sp4_v_b_14')
// (7, 6, 'sp4_v_b_3')
// (8, 1, 'sp4_r_v_b_36')
// (8, 2, 'sp12_h_r_14')
// (8, 2, 'sp4_h_r_21')
// (8, 2, 'sp4_r_v_b_25')
// (8, 3, 'sp4_r_v_b_12')
// (8, 4, 'sp4_h_r_42')
// (8, 4, 'sp4_h_r_43')
// (8, 4, 'sp4_r_v_b_1')
// (8, 5, 'local_g3_3')
// (8, 5, 'local_g3_6')
// (8, 5, 'lutff_1/in_2')
// (8, 5, 'lutff_4/in_2')
// (8, 5, 'lutff_6/in_2')
// (8, 5, 'sp4_r_v_b_43')
// (8, 5, 'sp4_r_v_b_46')
// (8, 6, 'sp4_r_v_b_30')
// (8, 6, 'sp4_r_v_b_35')
// (8, 7, 'sp4_r_v_b_19')
// (8, 7, 'sp4_r_v_b_22')
// (8, 8, 'sp4_r_v_b_11')
// (8, 8, 'sp4_r_v_b_6')
// (9, 0, 'span4_vert_36')
// (9, 1, 'sp4_v_b_36')
// (9, 2, 'sp12_h_r_17')
// (9, 2, 'sp4_h_r_32')
// (9, 2, 'sp4_v_b_25')
// (9, 3, 'sp4_v_b_12')
// (9, 4, 'local_g0_1')
// (9, 4, 'lutff_5/in_2')
// (9, 4, 'sp4_h_l_42')
// (9, 4, 'sp4_h_l_43')
// (9, 4, 'sp4_h_r_10')
// (9, 4, 'sp4_v_b_1')
// (9, 4, 'sp4_v_t_43')
// (9, 4, 'sp4_v_t_46')
// (9, 5, 'local_g2_6')
// (9, 5, 'local_g3_6')
// (9, 5, 'lutff_1/in_3')
// (9, 5, 'lutff_4/in_2')
// (9, 5, 'lutff_5/in_2')
// (9, 5, 'sp4_v_b_43')
// (9, 5, 'sp4_v_b_46')
// (9, 6, 'sp4_v_b_30')
// (9, 6, 'sp4_v_b_35')
// (9, 7, 'sp4_v_b_19')
// (9, 7, 'sp4_v_b_22')
// (9, 8, 'sp4_v_b_11')
// (9, 8, 'sp4_v_b_6')
// (10, 2, 'sp12_h_r_18')
// (10, 2, 'sp4_h_r_45')
// (10, 3, 'sp4_r_v_b_36')
// (10, 4, 'sp4_h_r_23')
// (10, 4, 'sp4_r_v_b_25')
// (10, 5, 'sp4_r_v_b_12')
// (10, 6, 'sp4_r_v_b_1')
// (11, 2, 'sp12_h_r_21')
// (11, 2, 'sp4_h_l_45')
// (11, 2, 'sp4_v_t_36')
// (11, 3, 'sp4_v_b_36')
// (11, 4, 'local_g2_2')
// (11, 4, 'lutff_2/in_2')
// (11, 4, 'lutff_6/in_2')
// (11, 4, 'sp4_h_r_34')
// (11, 4, 'sp4_v_b_25')
// (11, 5, 'local_g0_4')
// (11, 5, 'local_g1_4')
// (11, 5, 'lutff_0/in_2')
// (11, 5, 'lutff_1/in_2')
// (11, 5, 'lutff_3/in_2')
// (11, 5, 'sp4_v_b_12')
// (11, 6, 'sp4_v_b_1')
// (12, 2, 'sp12_h_r_22')
// (12, 4, 'sp4_h_r_47')
// (13, 2, 'span12_horz_22')
// (13, 4, 'span4_horz_47')

wire n42;
// (1, 2, 'sp4_h_r_7')
// (2, 2, 'local_g0_2')
// (2, 2, 'lutff_4/in_0')
// (2, 2, 'lutff_6/in_2')
// (2, 2, 'sp4_h_r_18')
// (3, 1, 'neigh_op_tnr_5')
// (3, 2, 'neigh_op_rgt_5')
// (3, 2, 'sp4_h_r_31')
// (3, 3, 'neigh_op_bnr_5')
// (4, 1, 'neigh_op_top_5')
// (4, 2, 'local_g2_5')
// (4, 2, 'lutff_1/in_0')
// (4, 2, 'lutff_5/out')
// (4, 2, 'sp4_h_r_42')
// (4, 3, 'neigh_op_bot_5')
// (5, 1, 'neigh_op_tnl_5')
// (5, 2, 'neigh_op_lft_5')
// (5, 2, 'sp4_h_l_42')
// (5, 3, 'neigh_op_bnl_5')

wire n43;
// (1, 3, 'neigh_op_tnr_1')
// (1, 4, 'neigh_op_rgt_1')
// (1, 5, 'neigh_op_bnr_1')
// (2, 3, 'neigh_op_top_1')
// (2, 4, 'local_g1_1')
// (2, 4, 'lutff_1/out')
// (2, 4, 'lutff_3/in_3')
// (2, 5, 'neigh_op_bot_1')
// (3, 3, 'neigh_op_tnl_1')
// (3, 4, 'neigh_op_lft_1')
// (3, 5, 'neigh_op_bnl_1')

wire n44;
// (1, 3, 'neigh_op_tnr_2')
// (1, 4, 'neigh_op_rgt_2')
// (1, 4, 'sp4_r_v_b_36')
// (1, 5, 'neigh_op_bnr_2')
// (1, 5, 'sp4_r_v_b_25')
// (1, 6, 'sp4_r_v_b_12')
// (1, 7, 'sp4_r_v_b_1')
// (2, 3, 'neigh_op_top_2')
// (2, 3, 'sp4_v_t_36')
// (2, 4, 'lutff_2/out')
// (2, 4, 'sp4_v_b_36')
// (2, 5, 'neigh_op_bot_2')
// (2, 5, 'sp4_v_b_25')
// (2, 6, 'local_g0_4')
// (2, 6, 'lutff_0/in_2')
// (2, 6, 'sp4_v_b_12')
// (2, 7, 'sp4_v_b_1')
// (3, 3, 'neigh_op_tnl_2')
// (3, 4, 'neigh_op_lft_2')
// (3, 5, 'neigh_op_bnl_2')

wire n45;
// (1, 3, 'neigh_op_tnr_3')
// (1, 4, 'neigh_op_rgt_3')
// (1, 5, 'neigh_op_bnr_3')
// (2, 3, 'neigh_op_top_3')
// (2, 4, 'lutff_3/out')
// (2, 4, 'sp4_h_r_6')
// (2, 5, 'neigh_op_bot_3')
// (3, 3, 'neigh_op_tnl_3')
// (3, 4, 'neigh_op_lft_3')
// (3, 4, 'sp4_h_r_19')
// (3, 5, 'neigh_op_bnl_3')
// (4, 4, 'sp4_h_r_30')
// (5, 4, 'sp4_h_r_43')
// (6, 4, 'sp4_h_l_43')
// (6, 4, 'sp4_h_r_9')
// (7, 4, 'local_g0_4')
// (7, 4, 'lutff_6/in_2')
// (7, 4, 'sp4_h_r_20')
// (8, 4, 'sp4_h_r_33')
// (9, 4, 'sp4_h_r_44')
// (10, 4, 'sp4_h_l_44')

wire n46;
// (1, 3, 'sp12_h_r_1')
// (2, 3, 'sp12_h_r_2')
// (3, 3, 'sp12_h_r_5')
// (4, 3, 'sp12_h_r_6')
// (5, 2, 'neigh_op_tnr_1')
// (5, 3, 'neigh_op_rgt_1')
// (5, 3, 'sp12_h_r_9')
// (5, 4, 'neigh_op_bnr_1')
// (6, 2, 'neigh_op_top_1')
// (6, 3, 'lutff_1/out')
// (6, 3, 'sp12_h_r_10')
// (6, 4, 'neigh_op_bot_1')
// (7, 2, 'neigh_op_tnl_1')
// (7, 3, 'neigh_op_lft_1')
// (7, 3, 'sp12_h_r_13')
// (7, 4, 'local_g2_1')
// (7, 4, 'lutff_5/in_0')
// (7, 4, 'neigh_op_bnl_1')
// (8, 3, 'local_g1_6')
// (8, 3, 'lutff_4/in_1')
// (8, 3, 'sp12_h_r_14')
// (9, 3, 'sp12_h_r_17')
// (10, 3, 'sp12_h_r_18')
// (11, 3, 'sp12_h_r_21')
// (12, 3, 'sp12_h_r_22')
// (13, 3, 'span12_horz_22')

wire n47;
// (1, 3, 'sp4_r_v_b_37')
// (1, 4, 'sp4_r_v_b_24')
// (1, 5, 'neigh_op_tnr_0')
// (1, 5, 'sp4_r_v_b_13')
// (1, 6, 'neigh_op_rgt_0')
// (1, 6, 'sp4_r_v_b_0')
// (1, 7, 'neigh_op_bnr_0')
// (1, 7, 'sp4_r_v_b_38')
// (1, 8, 'local_g1_3')
// (1, 8, 'lutff_global/cen')
// (1, 8, 'sp4_r_v_b_27')
// (1, 9, 'sp4_r_v_b_14')
// (1, 10, 'sp4_r_v_b_3')
// (2, 2, 'sp4_v_t_37')
// (2, 3, 'sp4_v_b_37')
// (2, 4, 'sp4_v_b_24')
// (2, 5, 'neigh_op_top_0')
// (2, 5, 'sp4_v_b_13')
// (2, 6, 'lutff_0/out')
// (2, 6, 'sp4_v_b_0')
// (2, 6, 'sp4_v_t_38')
// (2, 7, 'neigh_op_bot_0')
// (2, 7, 'sp4_v_b_38')
// (2, 8, 'sp4_v_b_27')
// (2, 9, 'sp4_v_b_14')
// (2, 10, 'sp4_v_b_3')
// (3, 5, 'neigh_op_tnl_0')
// (3, 6, 'neigh_op_lft_0')
// (3, 7, 'neigh_op_bnl_0')

reg n48 = 0;
// (1, 4, 'neigh_op_tnr_2')
// (1, 5, 'neigh_op_rgt_2')
// (1, 5, 'sp4_r_v_b_36')
// (1, 6, 'neigh_op_bnr_2')
// (1, 6, 'sp4_r_v_b_25')
// (1, 7, 'sp4_r_v_b_12')
// (1, 8, 'sp4_r_v_b_1')
// (2, 4, 'neigh_op_top_2')
// (2, 4, 'sp4_v_t_36')
// (2, 5, 'local_g0_2')
// (2, 5, 'lutff_2/in_2')
// (2, 5, 'lutff_2/out')
// (2, 5, 'sp4_v_b_36')
// (2, 6, 'local_g1_2')
// (2, 6, 'lutff_1/in_0')
// (2, 6, 'neigh_op_bot_2')
// (2, 6, 'sp4_v_b_25')
// (2, 7, 'local_g1_4')
// (2, 7, 'lutff_7/in_2')
// (2, 7, 'sp4_v_b_12')
// (2, 8, 'sp4_v_b_1')
// (3, 4, 'neigh_op_tnl_2')
// (3, 5, 'neigh_op_lft_2')
// (3, 6, 'neigh_op_bnl_2')

reg n49 = 0;
// (1, 4, 'neigh_op_tnr_3')
// (1, 5, 'neigh_op_rgt_3')
// (1, 5, 'sp4_r_v_b_38')
// (1, 6, 'neigh_op_bnr_3')
// (1, 6, 'sp4_r_v_b_27')
// (1, 7, 'sp4_r_v_b_14')
// (1, 8, 'sp4_r_v_b_3')
// (2, 4, 'neigh_op_top_3')
// (2, 4, 'sp4_v_t_38')
// (2, 5, 'local_g0_3')
// (2, 5, 'lutff_3/in_2')
// (2, 5, 'lutff_3/out')
// (2, 5, 'sp4_v_b_38')
// (2, 6, 'local_g0_3')
// (2, 6, 'lutff_1/in_2')
// (2, 6, 'neigh_op_bot_3')
// (2, 6, 'sp4_v_b_27')
// (2, 7, 'local_g1_6')
// (2, 7, 'lutff_4/in_1')
// (2, 7, 'lutff_7/in_0')
// (2, 7, 'sp4_v_b_14')
// (2, 8, 'sp4_v_b_3')
// (3, 4, 'neigh_op_tnl_3')
// (3, 5, 'neigh_op_lft_3')
// (3, 6, 'neigh_op_bnl_3')

reg n50 = 0;
// (1, 4, 'neigh_op_tnr_4')
// (1, 5, 'neigh_op_rgt_4')
// (1, 6, 'neigh_op_bnr_4')
// (2, 4, 'local_g1_4')
// (2, 4, 'lutff_2/in_3')
// (2, 4, 'lutff_3/in_0')
// (2, 4, 'neigh_op_top_4')
// (2, 5, 'local_g0_4')
// (2, 5, 'lutff_4/in_2')
// (2, 5, 'lutff_4/out')
// (2, 5, 'sp12_h_r_0')
// (2, 5, 'sp4_h_r_8')
// (2, 6, 'neigh_op_bot_4')
// (3, 4, 'neigh_op_tnl_4')
// (3, 5, 'neigh_op_lft_4')
// (3, 5, 'sp12_h_r_3')
// (3, 5, 'sp4_h_r_21')
// (3, 5, 'sp4_h_r_3')
// (3, 6, 'neigh_op_bnl_4')
// (4, 2, 'sp4_r_v_b_40')
// (4, 3, 'sp4_r_v_b_29')
// (4, 4, 'sp4_r_v_b_16')
// (4, 5, 'sp12_h_r_4')
// (4, 5, 'sp4_h_r_14')
// (4, 5, 'sp4_h_r_32')
// (4, 5, 'sp4_r_v_b_5')
// (5, 1, 'sp4_v_t_40')
// (5, 2, 'sp4_r_v_b_39')
// (5, 2, 'sp4_v_b_40')
// (5, 3, 'sp4_r_v_b_26')
// (5, 3, 'sp4_v_b_29')
// (5, 4, 'local_g0_0')
// (5, 4, 'lutff_5/in_1')
// (5, 4, 'sp4_r_v_b_15')
// (5, 4, 'sp4_v_b_16')
// (5, 5, 'sp12_h_r_7')
// (5, 5, 'sp4_h_r_27')
// (5, 5, 'sp4_h_r_45')
// (5, 5, 'sp4_h_r_5')
// (5, 5, 'sp4_r_v_b_2')
// (5, 5, 'sp4_v_b_5')
// (6, 1, 'sp4_v_t_39')
// (6, 2, 'sp4_r_v_b_38')
// (6, 2, 'sp4_v_b_39')
// (6, 3, 'sp4_r_v_b_27')
// (6, 3, 'sp4_v_b_26')
// (6, 4, 'local_g0_7')
// (6, 4, 'local_g2_6')
// (6, 4, 'lutff_2/in_1')
// (6, 4, 'lutff_4/in_3')
// (6, 4, 'lutff_5/in_1')
// (6, 4, 'sp4_r_v_b_14')
// (6, 4, 'sp4_v_b_15')
// (6, 5, 'local_g0_0')
// (6, 5, 'local_g2_6')
// (6, 5, 'lutff_2/in_0')
// (6, 5, 'lutff_4/in_2')
// (6, 5, 'lutff_5/in_3')
// (6, 5, 'sp12_h_r_8')
// (6, 5, 'sp4_h_l_45')
// (6, 5, 'sp4_h_r_16')
// (6, 5, 'sp4_h_r_38')
// (6, 5, 'sp4_r_v_b_3')
// (6, 5, 'sp4_v_b_2')
// (7, 1, 'sp4_v_t_38')
// (7, 2, 'sp4_v_b_38')
// (7, 3, 'sp4_v_b_27')
// (7, 4, 'sp4_v_b_14')
// (7, 5, 'sp12_h_r_11')
// (7, 5, 'sp4_h_l_38')
// (7, 5, 'sp4_h_r_29')
// (7, 5, 'sp4_v_b_3')
// (8, 5, 'sp12_h_r_12')
// (8, 5, 'sp4_h_r_40')
// (9, 5, 'sp12_h_r_15')
// (9, 5, 'sp4_h_l_40')
// (10, 5, 'sp12_h_r_16')
// (11, 5, 'sp12_h_r_19')
// (12, 5, 'sp12_h_r_20')
// (13, 5, 'span12_horz_20')

reg n51 = 0;
// (1, 4, 'neigh_op_tnr_5')
// (1, 5, 'neigh_op_rgt_5')
// (1, 5, 'sp12_h_r_1')
// (1, 6, 'neigh_op_bnr_5')
// (2, 4, 'local_g0_5')
// (2, 4, 'lutff_1/in_2')
// (2, 4, 'neigh_op_top_5')
// (2, 5, 'local_g0_5')
// (2, 5, 'lutff_5/in_2')
// (2, 5, 'lutff_5/out')
// (2, 5, 'sp12_h_r_2')
// (2, 5, 'sp4_h_r_10')
// (2, 6, 'neigh_op_bot_5')
// (3, 4, 'neigh_op_tnl_5')
// (3, 5, 'neigh_op_lft_5')
// (3, 5, 'sp12_h_r_5')
// (3, 5, 'sp4_h_r_23')
// (3, 6, 'neigh_op_bnl_5')
// (4, 2, 'sp4_r_v_b_44')
// (4, 3, 'sp4_r_v_b_33')
// (4, 4, 'sp4_r_v_b_20')
// (4, 5, 'sp12_h_r_6')
// (4, 5, 'sp4_h_r_34')
// (4, 5, 'sp4_r_v_b_9')
// (5, 1, 'sp4_v_t_44')
// (5, 2, 'sp4_r_v_b_41')
// (5, 2, 'sp4_v_b_44')
// (5, 3, 'sp4_r_v_b_28')
// (5, 3, 'sp4_v_b_33')
// (5, 4, 'local_g0_4')
// (5, 4, 'local_g1_4')
// (5, 4, 'lutff_2/in_3')
// (5, 4, 'lutff_5/in_3')
// (5, 4, 'sp4_r_v_b_17')
// (5, 4, 'sp4_v_b_20')
// (5, 5, 'sp12_h_r_9')
// (5, 5, 'sp4_h_r_4')
// (5, 5, 'sp4_h_r_47')
// (5, 5, 'sp4_r_v_b_4')
// (5, 5, 'sp4_v_b_9')
// (6, 1, 'sp4_v_t_41')
// (6, 2, 'sp4_v_b_41')
// (6, 3, 'sp4_v_b_28')
// (6, 4, 'local_g0_1')
// (6, 4, 'local_g1_1')
// (6, 4, 'lutff_0/in_1')
// (6, 4, 'lutff_4/in_2')
// (6, 4, 'sp4_v_b_17')
// (6, 5, 'local_g0_1')
// (6, 5, 'local_g0_2')
// (6, 5, 'lutff_2/in_1')
// (6, 5, 'lutff_4/in_1')
// (6, 5, 'lutff_5/in_1')
// (6, 5, 'sp12_h_r_10')
// (6, 5, 'sp4_h_l_47')
// (6, 5, 'sp4_h_r_17')
// (6, 5, 'sp4_v_b_4')
// (7, 5, 'sp12_h_r_13')
// (7, 5, 'sp4_h_r_28')
// (8, 5, 'sp12_h_r_14')
// (8, 5, 'sp4_h_r_41')
// (9, 5, 'sp12_h_r_17')
// (9, 5, 'sp4_h_l_41')
// (10, 5, 'sp12_h_r_18')
// (11, 5, 'sp12_h_r_21')
// (12, 5, 'sp12_h_r_22')
// (13, 5, 'span12_horz_22')

reg n52 = 0;
// (1, 4, 'neigh_op_tnr_6')
// (1, 5, 'neigh_op_rgt_6')
// (1, 5, 'sp4_h_r_0')
// (1, 5, 'sp4_h_r_1')
// (1, 6, 'neigh_op_bnr_6')
// (2, 4, 'local_g1_6')
// (2, 4, 'lutff_3/in_2')
// (2, 4, 'neigh_op_top_6')
// (2, 5, 'local_g0_6')
// (2, 5, 'lutff_6/in_2')
// (2, 5, 'lutff_6/out')
// (2, 5, 'sp4_h_r_12')
// (2, 5, 'sp4_h_r_13')
// (2, 5, 'sp4_r_v_b_45')
// (2, 6, 'neigh_op_bot_6')
// (2, 6, 'sp4_r_v_b_32')
// (2, 7, 'sp4_r_v_b_21')
// (2, 8, 'sp4_r_v_b_8')
// (3, 4, 'neigh_op_tnl_6')
// (3, 4, 'sp4_h_r_1')
// (3, 4, 'sp4_v_t_45')
// (3, 5, 'neigh_op_lft_6')
// (3, 5, 'sp4_h_r_24')
// (3, 5, 'sp4_h_r_25')
// (3, 5, 'sp4_v_b_45')
// (3, 6, 'neigh_op_bnl_6')
// (3, 6, 'sp4_v_b_32')
// (3, 7, 'sp4_v_b_21')
// (3, 8, 'sp4_v_b_8')
// (4, 2, 'sp4_r_v_b_42')
// (4, 3, 'sp4_r_v_b_31')
// (4, 4, 'sp4_h_r_12')
// (4, 4, 'sp4_r_v_b_18')
// (4, 5, 'sp4_h_r_36')
// (4, 5, 'sp4_h_r_37')
// (4, 5, 'sp4_r_v_b_7')
// (5, 1, 'sp4_v_t_42')
// (5, 2, 'sp4_v_b_42')
// (5, 3, 'sp4_v_b_31')
// (5, 4, 'local_g0_2')
// (5, 4, 'local_g1_2')
// (5, 4, 'lutff_2/in_2')
// (5, 4, 'lutff_5/in_0')
// (5, 4, 'sp4_h_r_25')
// (5, 4, 'sp4_v_b_18')
// (5, 5, 'sp4_h_l_36')
// (5, 5, 'sp4_h_l_37')
// (5, 5, 'sp4_h_r_0')
// (5, 5, 'sp4_v_b_7')
// (6, 4, 'local_g2_4')
// (6, 4, 'lutff_0/in_2')
// (6, 4, 'sp4_h_r_36')
// (6, 5, 'local_g0_5')
// (6, 5, 'lutff_3/in_0')
// (6, 5, 'lutff_5/in_0')
// (6, 5, 'lutff_6/in_3')
// (6, 5, 'sp4_h_r_13')
// (7, 4, 'sp4_h_l_36')
// (7, 5, 'sp4_h_r_24')
// (8, 5, 'sp4_h_r_37')
// (9, 5, 'sp4_h_l_37')

wire n53;
// (1, 5, 'neigh_op_tnr_1')
// (1, 6, 'neigh_op_rgt_1')
// (1, 7, 'neigh_op_bnr_1')
// (2, 5, 'neigh_op_top_1')
// (2, 6, 'local_g0_1')
// (2, 6, 'lutff_0/in_1')
// (2, 6, 'lutff_1/out')
// (2, 7, 'neigh_op_bot_1')
// (3, 5, 'neigh_op_tnl_1')
// (3, 6, 'neigh_op_lft_1')
// (3, 7, 'neigh_op_bnl_1')

wire n54;
// (1, 5, 'neigh_op_tnr_3')
// (1, 6, 'neigh_op_rgt_3')
// (1, 7, 'neigh_op_bnr_3')
// (2, 4, 'sp4_r_v_b_47')
// (2, 5, 'neigh_op_top_3')
// (2, 5, 'sp4_r_v_b_34')
// (2, 6, 'lutff_3/out')
// (2, 6, 'sp4_r_v_b_23')
// (2, 7, 'neigh_op_bot_3')
// (2, 7, 'sp4_r_v_b_10')
// (3, 3, 'sp4_v_t_47')
// (3, 4, 'sp4_v_b_47')
// (3, 5, 'neigh_op_tnl_3')
// (3, 5, 'sp4_v_b_34')
// (3, 6, 'neigh_op_lft_3')
// (3, 6, 'sp4_v_b_23')
// (3, 7, 'neigh_op_bnl_3')
// (3, 7, 'sp4_h_r_10')
// (3, 7, 'sp4_h_r_4')
// (3, 7, 'sp4_v_b_10')
// (4, 7, 'local_g1_1')
// (4, 7, 'lutff_6/in_2')
// (4, 7, 'lutff_7/in_3')
// (4, 7, 'sp4_h_r_17')
// (4, 7, 'sp4_h_r_23')
// (5, 7, 'local_g2_4')
// (5, 7, 'lutff_3/in_3')
// (5, 7, 'lutff_7/in_1')
// (5, 7, 'sp4_h_r_28')
// (5, 7, 'sp4_h_r_34')
// (6, 7, 'local_g2_1')
// (6, 7, 'local_g3_7')
// (6, 7, 'lutff_0/in_1')
// (6, 7, 'lutff_1/in_3')
// (6, 7, 'lutff_4/in_1')
// (6, 7, 'lutff_6/in_0')
// (6, 7, 'sp4_h_r_41')
// (6, 7, 'sp4_h_r_47')
// (7, 7, 'sp4_h_l_41')
// (7, 7, 'sp4_h_l_47')

reg n55 = 0;
// (1, 5, 'neigh_op_tnr_7')
// (1, 6, 'neigh_op_rgt_7')
// (1, 7, 'neigh_op_bnr_7')
// (2, 5, 'local_g0_7')
// (2, 5, 'lutff_1/in_2')
// (2, 5, 'neigh_op_top_7')
// (2, 6, 'local_g0_7')
// (2, 6, 'local_g1_7')
// (2, 6, 'lutff_1/in_3')
// (2, 6, 'lutff_7/in_2')
// (2, 6, 'lutff_7/out')
// (2, 7, 'local_g0_7')
// (2, 7, 'local_g1_7')
// (2, 7, 'lutff_0/in_3')
// (2, 7, 'lutff_4/in_3')
// (2, 7, 'lutff_7/in_1')
// (2, 7, 'neigh_op_bot_7')
// (3, 5, 'neigh_op_tnl_7')
// (3, 6, 'neigh_op_lft_7')
// (3, 7, 'neigh_op_bnl_7')

reg n56 = 0;
// (1, 5, 'sp12_h_r_0')
// (2, 5, 'sp12_h_r_3')
// (3, 5, 'sp12_h_r_4')
// (4, 5, 'sp12_h_r_7')
// (4, 5, 'sp4_h_r_5')
// (5, 5, 'sp12_h_r_8')
// (5, 5, 'sp4_h_r_16')
// (6, 5, 'sp12_h_r_11')
// (6, 5, 'sp4_h_r_29')
// (7, 5, 'local_g2_0')
// (7, 5, 'lutff_6/in_0')
// (7, 5, 'sp12_h_r_12')
// (7, 5, 'sp4_h_r_40')
// (8, 5, 'sp12_h_r_15')
// (8, 5, 'sp4_h_l_40')
// (9, 5, 'sp12_h_r_16')
// (10, 4, 'neigh_op_tnr_6')
// (10, 5, 'neigh_op_rgt_6')
// (10, 5, 'sp12_h_r_19')
// (10, 6, 'neigh_op_bnr_6')
// (11, 4, 'local_g1_6')
// (11, 4, 'lutff_6/in_3')
// (11, 4, 'neigh_op_top_6')
// (11, 5, 'lutff_6/out')
// (11, 5, 'sp12_h_r_20')
// (11, 6, 'neigh_op_bot_6')
// (12, 4, 'neigh_op_tnl_6')
// (12, 5, 'neigh_op_lft_6')
// (12, 5, 'sp12_h_r_23')
// (12, 6, 'neigh_op_bnl_6')
// (13, 5, 'span12_horz_23')

wire n57;
// (1, 5, 'sp4_r_v_b_40')
// (1, 6, 'neigh_op_tnr_0')
// (1, 6, 'sp4_r_v_b_29')
// (1, 7, 'neigh_op_rgt_0')
// (1, 7, 'sp4_r_v_b_16')
// (1, 8, 'neigh_op_bnr_0')
// (1, 8, 'sp4_r_v_b_5')
// (2, 4, 'sp4_v_t_40')
// (2, 5, 'sp4_v_b_40')
// (2, 6, 'neigh_op_top_0')
// (2, 6, 'sp4_v_b_29')
// (2, 7, 'local_g0_0')
// (2, 7, 'lutff_0/out')
// (2, 7, 'lutff_6/in_0')
// (2, 7, 'sp4_v_b_16')
// (2, 8, 'local_g1_5')
// (2, 8, 'lutff_7/in_3')
// (2, 8, 'neigh_op_bot_0')
// (2, 8, 'sp4_v_b_5')
// (3, 6, 'neigh_op_tnl_0')
// (3, 7, 'neigh_op_lft_0')
// (3, 8, 'neigh_op_bnl_0')

reg n58 = 0;
// (1, 5, 'sp4_r_v_b_44')
// (1, 6, 'sp4_r_v_b_33')
// (1, 7, 'sp4_r_v_b_20')
// (1, 8, 'sp4_r_v_b_9')
// (2, 4, 'sp4_h_r_3')
// (2, 4, 'sp4_v_t_44')
// (2, 5, 'sp4_v_b_44')
// (2, 6, 'sp4_v_b_33')
// (2, 7, 'local_g0_4')
// (2, 7, 'lutff_global/s_r')
// (2, 7, 'sp4_v_b_20')
// (2, 8, 'sp4_v_b_9')
// (3, 4, 'sp4_h_r_14')
// (4, 1, 'neigh_op_tnr_5')
// (4, 2, 'local_g3_5')
// (4, 2, 'lutff_2/in_2')
// (4, 2, 'lutff_4/in_0')
// (4, 2, 'neigh_op_rgt_5')
// (4, 3, 'local_g0_5')
// (4, 3, 'lutff_4/in_1')
// (4, 3, 'neigh_op_bnr_5')
// (4, 4, 'sp4_h_r_27')
// (5, 1, 'neigh_op_top_5')
// (5, 1, 'sp4_r_v_b_38')
// (5, 2, 'local_g0_5')
// (5, 2, 'lutff_4/in_1')
// (5, 2, 'lutff_5/in_2')
// (5, 2, 'lutff_5/out')
// (5, 2, 'sp4_r_v_b_27')
// (5, 3, 'neigh_op_bot_5')
// (5, 3, 'sp4_r_v_b_14')
// (5, 4, 'sp4_h_r_38')
// (5, 4, 'sp4_r_v_b_3')
// (6, 0, 'span4_vert_38')
// (6, 1, 'neigh_op_tnl_5')
// (6, 1, 'sp4_v_b_38')
// (6, 2, 'neigh_op_lft_5')
// (6, 2, 'sp4_v_b_27')
// (6, 3, 'neigh_op_bnl_5')
// (6, 3, 'sp4_v_b_14')
// (6, 4, 'sp4_h_l_38')
// (6, 4, 'sp4_v_b_3')

reg n59 = 0;
// (1, 6, 'neigh_op_tnr_4')
// (1, 6, 'sp4_r_v_b_37')
// (1, 7, 'neigh_op_rgt_4')
// (1, 7, 'sp4_r_v_b_24')
// (1, 8, 'neigh_op_bnr_4')
// (1, 8, 'sp4_r_v_b_13')
// (1, 9, 'sp4_r_v_b_0')
// (1, 10, 'sp4_r_v_b_37')
// (1, 11, 'sp4_r_v_b_24')
// (1, 12, 'sp4_r_v_b_13')
// (1, 13, 'sp4_r_v_b_0')
// (2, 0, 'span12_vert_20')
// (2, 1, 'sp12_v_b_20')
// (2, 2, 'sp12_v_b_19')
// (2, 3, 'sp12_v_b_16')
// (2, 4, 'sp12_v_b_15')
// (2, 5, 'sp12_v_b_12')
// (2, 5, 'sp4_v_t_37')
// (2, 6, 'neigh_op_top_4')
// (2, 6, 'sp12_v_b_11')
// (2, 6, 'sp4_v_b_37')
// (2, 7, 'lutff_4/out')
// (2, 7, 'sp12_v_b_8')
// (2, 7, 'sp4_v_b_24')
// (2, 8, 'neigh_op_bot_4')
// (2, 8, 'sp12_v_b_7')
// (2, 8, 'sp4_v_b_13')
// (2, 9, 'sp12_v_b_4')
// (2, 9, 'sp4_h_r_6')
// (2, 9, 'sp4_v_b_0')
// (2, 9, 'sp4_v_t_37')
// (2, 10, 'sp12_v_b_3')
// (2, 10, 'sp4_v_b_37')
// (2, 11, 'sp12_h_r_0')
// (2, 11, 'sp12_v_b_0')
// (2, 11, 'sp4_v_b_24')
// (2, 12, 'sp4_v_b_13')
// (2, 13, 'local_g0_0')
// (2, 13, 'lutff_0/in_2')
// (2, 13, 'sp4_h_r_0')
// (2, 13, 'sp4_v_b_0')
// (3, 6, 'neigh_op_tnl_4')
// (3, 7, 'neigh_op_lft_4')
// (3, 8, 'neigh_op_bnl_4')
// (3, 9, 'sp4_h_r_19')
// (3, 11, 'sp12_h_r_3')
// (3, 11, 'sp4_h_r_3')
// (3, 13, 'sp4_h_r_13')
// (4, 9, 'sp4_h_r_30')
// (4, 11, 'sp12_h_r_4')
// (4, 11, 'sp4_h_r_14')
// (4, 13, 'local_g2_0')
// (4, 13, 'local_g3_0')
// (4, 13, 'lutff_0/in_3')
// (4, 13, 'lutff_5/in_3')
// (4, 13, 'sp4_h_r_24')
// (5, 9, 'local_g2_3')
// (5, 9, 'lutff_2/in_3')
// (5, 9, 'sp4_h_r_43')
// (5, 10, 'sp4_r_v_b_37')
// (5, 11, 'local_g1_0')
// (5, 11, 'lutff_6/in_3')
// (5, 11, 'sp12_h_r_7')
// (5, 11, 'sp4_h_r_27')
// (5, 11, 'sp4_r_v_b_24')
// (5, 12, 'local_g2_5')
// (5, 12, 'lutff_1/in_2')
// (5, 12, 'sp4_r_v_b_13')
// (5, 13, 'local_g2_5')
// (5, 13, 'local_g3_5')
// (5, 13, 'lutff_0/in_2')
// (5, 13, 'lutff_1/in_3')
// (5, 13, 'lutff_7/in_2')
// (5, 13, 'sp4_h_r_37')
// (5, 13, 'sp4_r_v_b_0')
// (5, 14, 'local_g2_5')
// (5, 14, 'lutff_4/in_3')
// (5, 14, 'sp4_r_v_b_37')
// (5, 15, 'sp4_r_v_b_24')
// (5, 16, 'sp4_r_v_b_13')
// (6, 9, 'sp4_h_l_43')
// (6, 9, 'sp4_h_r_5')
// (6, 9, 'sp4_v_t_37')
// (6, 10, 'sp4_v_b_37')
// (6, 11, 'sp12_h_r_8')
// (6, 11, 'sp4_h_r_38')
// (6, 11, 'sp4_v_b_24')
// (6, 12, 'local_g1_5')
// (6, 12, 'lutff_0/in_2')
// (6, 12, 'lutff_1/in_3')
// (6, 12, 'lutff_2/in_2')
// (6, 12, 'sp4_r_v_b_45')
// (6, 12, 'sp4_v_b_13')
// (6, 13, 'local_g1_0')
// (6, 13, 'lutff_2/in_3')
// (6, 13, 'sp4_h_l_37')
// (6, 13, 'sp4_h_r_5')
// (6, 13, 'sp4_r_v_b_32')
// (6, 13, 'sp4_v_b_0')
// (6, 13, 'sp4_v_t_37')
// (6, 14, 'local_g2_5')
// (6, 14, 'local_g3_5')
// (6, 14, 'lutff_0/in_3')
// (6, 14, 'lutff_1/in_2')
// (6, 14, 'lutff_3/in_2')
// (6, 14, 'lutff_5/in_3')
// (6, 14, 'sp4_r_v_b_21')
// (6, 14, 'sp4_v_b_37')
// (6, 15, 'local_g2_0')
// (6, 15, 'lutff_7/in_3')
// (6, 15, 'sp4_r_v_b_8')
// (6, 15, 'sp4_v_b_24')
// (6, 16, 'sp4_v_b_13')
// (6, 17, 'span4_vert_0')
// (7, 9, 'local_g0_0')
// (7, 9, 'lutff_2/in_2')
// (7, 9, 'sp4_h_r_16')
// (7, 11, 'local_g0_3')
// (7, 11, 'lutff_0/in_3')
// (7, 11, 'lutff_7/in_2')
// (7, 11, 'sp12_h_r_11')
// (7, 11, 'sp4_h_l_38')
// (7, 11, 'sp4_v_t_45')
// (7, 12, 'sp4_v_b_45')
// (7, 13, 'local_g0_0')
// (7, 13, 'local_g1_0')
// (7, 13, 'lutff_0/in_2')
// (7, 13, 'lutff_4/in_3')
// (7, 13, 'lutff_5/in_2')
// (7, 13, 'sp4_h_r_16')
// (7, 13, 'sp4_v_b_32')
// (7, 14, 'local_g0_5')
// (7, 14, 'lutff_0/in_3')
// (7, 14, 'lutff_3/in_2')
// (7, 14, 'sp4_v_b_21')
// (7, 15, 'local_g0_2')
// (7, 15, 'lutff_3/in_3')
// (7, 15, 'sp4_h_r_2')
// (7, 15, 'sp4_v_b_8')
// (8, 9, 'local_g2_5')
// (8, 9, 'local_g3_5')
// (8, 9, 'lutff_0/in_2')
// (8, 9, 'lutff_1/in_3')
// (8, 9, 'lutff_3/in_2')
// (8, 9, 'sp4_h_r_29')
// (8, 11, 'local_g0_4')
// (8, 11, 'lutff_7/in_3')
// (8, 11, 'sp12_h_r_12')
// (8, 13, 'local_g2_5')
// (8, 13, 'lutff_1/in_2')
// (8, 13, 'sp4_h_r_29')
// (8, 15, 'sp4_h_r_15')
// (9, 9, 'sp4_h_r_40')
// (9, 11, 'sp12_h_r_15')
// (9, 13, 'sp4_h_r_40')
// (9, 15, 'sp4_h_r_26')
// (10, 9, 'sp4_h_l_40')
// (10, 11, 'sp12_h_r_16')
// (10, 13, 'sp4_h_l_40')
// (10, 15, 'sp4_h_r_39')
// (11, 11, 'sp12_h_r_19')
// (11, 15, 'sp4_h_l_39')
// (12, 11, 'sp12_h_r_20')
// (13, 11, 'span12_horz_20')

reg n60 = 0;
// (1, 6, 'neigh_op_tnr_7')
// (1, 7, 'neigh_op_rgt_7')
// (1, 7, 'sp4_h_r_3')
// (1, 8, 'neigh_op_bnr_7')
// (2, 2, 'sp12_v_t_22')
// (2, 3, 'sp12_v_b_22')
// (2, 4, 'sp12_v_b_21')
// (2, 5, 'sp12_v_b_18')
// (2, 6, 'neigh_op_top_7')
// (2, 6, 'sp12_v_b_17')
// (2, 7, 'lutff_7/out')
// (2, 7, 'sp12_v_b_14')
// (2, 7, 'sp4_h_r_14')
// (2, 8, 'neigh_op_bot_7')
// (2, 8, 'sp12_v_b_13')
// (2, 9, 'sp12_v_b_10')
// (2, 10, 'sp12_v_b_9')
// (2, 11, 'sp12_v_b_6')
// (2, 12, 'sp12_v_b_5')
// (2, 13, 'local_g3_2')
// (2, 13, 'lutff_0/in_3')
// (2, 13, 'sp12_v_b_2')
// (2, 14, 'sp12_h_r_1')
// (2, 14, 'sp12_v_b_1')
// (3, 6, 'neigh_op_tnl_7')
// (3, 7, 'neigh_op_lft_7')
// (3, 7, 'sp4_h_r_27')
// (3, 8, 'neigh_op_bnl_7')
// (3, 11, 'sp4_r_v_b_42')
// (3, 12, 'sp4_r_v_b_31')
// (3, 13, 'sp4_r_v_b_18')
// (3, 14, 'sp12_h_r_2')
// (3, 14, 'sp4_r_v_b_7')
// (4, 7, 'sp4_h_r_38')
// (4, 8, 'sp4_r_v_b_45')
// (4, 9, 'sp4_r_v_b_32')
// (4, 10, 'sp4_r_v_b_21')
// (4, 10, 'sp4_v_t_42')
// (4, 11, 'sp4_r_v_b_8')
// (4, 11, 'sp4_v_b_42')
// (4, 12, 'sp4_r_v_b_46')
// (4, 12, 'sp4_v_b_31')
// (4, 13, 'local_g0_2')
// (4, 13, 'local_g1_2')
// (4, 13, 'lutff_0/in_2')
// (4, 13, 'lutff_5/in_2')
// (4, 13, 'sp4_r_v_b_35')
// (4, 13, 'sp4_v_b_18')
// (4, 14, 'sp12_h_r_5')
// (4, 14, 'sp4_h_r_2')
// (4, 14, 'sp4_r_v_b_22')
// (4, 14, 'sp4_v_b_7')
// (4, 15, 'sp4_r_v_b_11')
// (5, 7, 'sp4_h_l_38')
// (5, 7, 'sp4_v_t_45')
// (5, 8, 'sp4_v_b_45')
// (5, 9, 'local_g2_0')
// (5, 9, 'lutff_2/in_2')
// (5, 9, 'sp4_v_b_32')
// (5, 10, 'sp4_v_b_21')
// (5, 11, 'local_g0_0')
// (5, 11, 'lutff_6/in_2')
// (5, 11, 'sp4_r_v_b_44')
// (5, 11, 'sp4_v_b_8')
// (5, 11, 'sp4_v_t_46')
// (5, 12, 'local_g2_6')
// (5, 12, 'lutff_1/in_1')
// (5, 12, 'sp4_r_v_b_33')
// (5, 12, 'sp4_v_b_46')
// (5, 13, 'local_g2_3')
// (5, 13, 'local_g3_3')
// (5, 13, 'lutff_0/in_1')
// (5, 13, 'lutff_1/in_2')
// (5, 13, 'lutff_7/in_3')
// (5, 13, 'sp4_r_v_b_20')
// (5, 13, 'sp4_v_b_35')
// (5, 14, 'local_g0_6')
// (5, 14, 'lutff_4/in_2')
// (5, 14, 'sp12_h_r_6')
// (5, 14, 'sp4_h_r_15')
// (5, 14, 'sp4_r_v_b_9')
// (5, 14, 'sp4_v_b_22')
// (5, 15, 'sp4_h_r_5')
// (5, 15, 'sp4_v_b_11')
// (6, 10, 'sp4_v_t_44')
// (6, 11, 'sp4_v_b_44')
// (6, 12, 'local_g2_1')
// (6, 12, 'lutff_0/in_1')
// (6, 12, 'lutff_1/in_2')
// (6, 12, 'lutff_2/in_3')
// (6, 12, 'sp4_v_b_33')
// (6, 13, 'local_g0_4')
// (6, 13, 'lutff_2/in_2')
// (6, 13, 'sp4_v_b_20')
// (6, 14, 'local_g0_1')
// (6, 14, 'local_g1_1')
// (6, 14, 'lutff_0/in_2')
// (6, 14, 'lutff_1/in_1')
// (6, 14, 'lutff_3/in_3')
// (6, 14, 'lutff_5/in_2')
// (6, 14, 'sp12_h_r_9')
// (6, 14, 'sp4_h_r_26')
// (6, 14, 'sp4_h_r_4')
// (6, 14, 'sp4_v_b_9')
// (6, 15, 'local_g1_0')
// (6, 15, 'lutff_7/in_2')
// (6, 15, 'sp4_h_r_16')
// (7, 7, 'sp4_r_v_b_46')
// (7, 8, 'sp4_r_v_b_35')
// (7, 9, 'local_g3_6')
// (7, 9, 'lutff_2/in_1')
// (7, 9, 'sp4_r_v_b_22')
// (7, 10, 'sp4_r_v_b_11')
// (7, 11, 'local_g3_5')
// (7, 11, 'lutff_0/in_2')
// (7, 11, 'lutff_7/in_3')
// (7, 11, 'sp4_r_v_b_39')
// (7, 11, 'sp4_r_v_b_45')
// (7, 12, 'sp4_r_v_b_26')
// (7, 12, 'sp4_r_v_b_32')
// (7, 13, 'local_g2_7')
// (7, 13, 'local_g3_5')
// (7, 13, 'lutff_0/in_1')
// (7, 13, 'lutff_4/in_2')
// (7, 13, 'lutff_5/in_1')
// (7, 13, 'sp4_r_v_b_15')
// (7, 13, 'sp4_r_v_b_21')
// (7, 14, 'local_g0_2')
// (7, 14, 'lutff_0/in_2')
// (7, 14, 'lutff_3/in_3')
// (7, 14, 'sp12_h_r_10')
// (7, 14, 'sp4_h_r_17')
// (7, 14, 'sp4_h_r_39')
// (7, 14, 'sp4_r_v_b_2')
// (7, 14, 'sp4_r_v_b_8')
// (7, 15, 'local_g2_7')
// (7, 15, 'lutff_3/in_2')
// (7, 15, 'sp4_h_r_29')
// (7, 15, 'sp4_r_v_b_39')
// (7, 16, 'sp4_r_v_b_26')
// (8, 6, 'sp4_v_t_46')
// (8, 7, 'sp4_v_b_46')
// (8, 8, 'sp4_v_b_35')
// (8, 9, 'local_g0_6')
// (8, 9, 'local_g1_6')
// (8, 9, 'lutff_0/in_1')
// (8, 9, 'lutff_1/in_2')
// (8, 9, 'lutff_3/in_3')
// (8, 9, 'sp4_v_b_22')
// (8, 10, 'sp4_v_b_11')
// (8, 10, 'sp4_v_t_39')
// (8, 10, 'sp4_v_t_45')
// (8, 11, 'local_g2_5')
// (8, 11, 'lutff_7/in_2')
// (8, 11, 'sp4_v_b_39')
// (8, 11, 'sp4_v_b_45')
// (8, 12, 'sp4_v_b_26')
// (8, 12, 'sp4_v_b_32')
// (8, 13, 'local_g1_5')
// (8, 13, 'lutff_1/in_3')
// (8, 13, 'sp4_v_b_15')
// (8, 13, 'sp4_v_b_21')
// (8, 14, 'sp12_h_r_13')
// (8, 14, 'sp4_h_l_39')
// (8, 14, 'sp4_h_r_28')
// (8, 14, 'sp4_v_b_2')
// (8, 14, 'sp4_v_b_8')
// (8, 14, 'sp4_v_t_39')
// (8, 15, 'sp4_h_r_40')
// (8, 15, 'sp4_v_b_39')
// (8, 16, 'sp4_v_b_26')
// (8, 17, 'span4_vert_15')
// (9, 14, 'sp12_h_r_14')
// (9, 14, 'sp4_h_r_41')
// (9, 15, 'sp4_h_l_40')
// (10, 14, 'sp12_h_r_17')
// (10, 14, 'sp4_h_l_41')
// (11, 14, 'sp12_h_r_18')
// (12, 14, 'sp12_h_r_21')
// (13, 14, 'span12_horz_21')

reg n61 = 0;
// (1, 7, 'neigh_op_tnr_2')
// (1, 8, 'neigh_op_rgt_2')
// (1, 8, 'sp4_h_r_9')
// (1, 8, 'sp4_r_v_b_36')
// (1, 9, 'neigh_op_bnr_2')
// (1, 9, 'sp4_r_v_b_25')
// (1, 10, 'sp4_r_v_b_12')
// (1, 11, 'sp4_r_v_b_1')
// (2, 7, 'neigh_op_top_2')
// (2, 7, 'sp4_v_t_36')
// (2, 8, 'lutff_2/out')
// (2, 8, 'sp4_h_r_20')
// (2, 8, 'sp4_v_b_36')
// (2, 9, 'neigh_op_bot_2')
// (2, 9, 'sp4_v_b_25')
// (2, 10, 'local_g1_4')
// (2, 10, 'lutff_7/in_0')
// (2, 10, 'sp4_v_b_12')
// (2, 11, 'sp4_v_b_1')
// (3, 7, 'neigh_op_tnl_2')
// (3, 8, 'neigh_op_lft_2')
// (3, 8, 'sp4_h_r_33')
// (3, 9, 'neigh_op_bnl_2')
// (4, 8, 'local_g3_4')
// (4, 8, 'lutff_2/in_1')
// (4, 8, 'sp4_h_r_44')
// (5, 8, 'sp4_h_l_44')

reg n62 = 0;
// (1, 7, 'neigh_op_tnr_7')
// (1, 8, 'neigh_op_rgt_7')
// (1, 8, 'sp4_h_r_0')
// (1, 8, 'sp4_h_r_3')
// (1, 9, 'neigh_op_bnr_7')
// (2, 6, 'sp4_r_v_b_39')
// (2, 7, 'neigh_op_top_7')
// (2, 7, 'sp4_r_v_b_26')
// (2, 8, 'local_g1_7')
// (2, 8, 'lutff_2/in_2')
// (2, 8, 'lutff_7/out')
// (2, 8, 'sp4_h_r_13')
// (2, 8, 'sp4_h_r_14')
// (2, 8, 'sp4_r_v_b_15')
// (2, 8, 'sp4_r_v_b_47')
// (2, 9, 'local_g0_1')
// (2, 9, 'lutff_3/in_2')
// (2, 9, 'neigh_op_bot_7')
// (2, 9, 'sp4_r_v_b_2')
// (2, 9, 'sp4_r_v_b_34')
// (2, 10, 'sp4_r_v_b_23')
// (2, 11, 'sp4_r_v_b_10')
// (3, 5, 'sp4_v_t_39')
// (3, 6, 'sp4_v_b_39')
// (3, 7, 'neigh_op_tnl_7')
// (3, 7, 'sp4_v_b_26')
// (3, 7, 'sp4_v_t_47')
// (3, 8, 'neigh_op_lft_7')
// (3, 8, 'sp4_h_r_24')
// (3, 8, 'sp4_h_r_27')
// (3, 8, 'sp4_v_b_15')
// (3, 8, 'sp4_v_b_47')
// (3, 9, 'neigh_op_bnl_7')
// (3, 9, 'sp4_h_r_2')
// (3, 9, 'sp4_v_b_2')
// (3, 9, 'sp4_v_b_34')
// (3, 10, 'sp4_v_b_23')
// (3, 11, 'sp4_h_r_10')
// (3, 11, 'sp4_v_b_10')
// (4, 5, 'sp4_r_v_b_38')
// (4, 6, 'sp4_r_v_b_27')
// (4, 7, 'sp4_r_v_b_14')
// (4, 8, 'local_g1_3')
// (4, 8, 'lutff_2/in_0')
// (4, 8, 'sp4_h_r_37')
// (4, 8, 'sp4_h_r_38')
// (4, 8, 'sp4_r_v_b_3')
// (4, 9, 'local_g0_7')
// (4, 9, 'local_g2_6')
// (4, 9, 'lutff_2/in_2')
// (4, 9, 'lutff_3/in_2')
// (4, 9, 'lutff_4/in_2')
// (4, 9, 'sp4_h_r_15')
// (4, 9, 'sp4_r_v_b_38')
// (4, 9, 'sp4_r_v_b_40')
// (4, 9, 'sp4_r_v_b_43')
// (4, 10, 'local_g1_5')
// (4, 10, 'local_g1_6')
// (4, 10, 'lutff_2/in_0')
// (4, 10, 'lutff_3/in_2')
// (4, 10, 'lutff_4/in_2')
// (4, 10, 'lutff_5/in_1')
// (4, 10, 'sp4_r_v_b_27')
// (4, 10, 'sp4_r_v_b_29')
// (4, 10, 'sp4_r_v_b_30')
// (4, 11, 'local_g0_7')
// (4, 11, 'lutff_3/in_2')
// (4, 11, 'lutff_5/in_2')
// (4, 11, 'sp4_h_r_23')
// (4, 11, 'sp4_r_v_b_14')
// (4, 11, 'sp4_r_v_b_16')
// (4, 11, 'sp4_r_v_b_19')
// (4, 12, 'sp4_r_v_b_3')
// (4, 12, 'sp4_r_v_b_5')
// (4, 12, 'sp4_r_v_b_6')
// (5, 4, 'sp4_v_t_38')
// (5, 5, 'sp4_v_b_38')
// (5, 6, 'sp4_v_b_27')
// (5, 7, 'sp4_v_b_14')
// (5, 8, 'sp4_h_l_37')
// (5, 8, 'sp4_h_l_38')
// (5, 8, 'sp4_h_r_8')
// (5, 8, 'sp4_v_b_3')
// (5, 8, 'sp4_v_t_38')
// (5, 8, 'sp4_v_t_40')
// (5, 8, 'sp4_v_t_43')
// (5, 9, 'local_g3_6')
// (5, 9, 'lutff_5/in_0')
// (5, 9, 'sp4_h_r_26')
// (5, 9, 'sp4_v_b_38')
// (5, 9, 'sp4_v_b_40')
// (5, 9, 'sp4_v_b_43')
// (5, 10, 'sp4_v_b_27')
// (5, 10, 'sp4_v_b_29')
// (5, 10, 'sp4_v_b_30')
// (5, 11, 'sp4_h_r_34')
// (5, 11, 'sp4_v_b_14')
// (5, 11, 'sp4_v_b_16')
// (5, 11, 'sp4_v_b_19')
// (5, 12, 'sp4_v_b_3')
// (5, 12, 'sp4_v_b_5')
// (5, 12, 'sp4_v_b_6')
// (6, 8, 'local_g3_1')
// (6, 8, 'lutff_3/in_1')
// (6, 8, 'sp4_h_r_21')
// (6, 8, 'sp4_r_v_b_41')
// (6, 8, 'sp4_r_v_b_47')
// (6, 9, 'local_g2_7')
// (6, 9, 'local_g3_7')
// (6, 9, 'lutff_4/in_2')
// (6, 9, 'lutff_5/in_2')
// (6, 9, 'lutff_7/in_2')
// (6, 9, 'sp4_h_r_39')
// (6, 9, 'sp4_r_v_b_28')
// (6, 9, 'sp4_r_v_b_34')
// (6, 10, 'local_g2_7')
// (6, 10, 'local_g3_1')
// (6, 10, 'lutff_1/in_2')
// (6, 10, 'lutff_4/in_2')
// (6, 10, 'lutff_6/in_1')
// (6, 10, 'lutff_7/in_2')
// (6, 10, 'sp4_r_v_b_17')
// (6, 10, 'sp4_r_v_b_23')
// (6, 10, 'sp4_r_v_b_39')
// (6, 11, 'local_g2_2')
// (6, 11, 'local_g2_7')
// (6, 11, 'lutff_2/in_2')
// (6, 11, 'lutff_4/in_2')
// (6, 11, 'lutff_6/in_2')
// (6, 11, 'lutff_7/in_0')
// (6, 11, 'sp4_h_r_47')
// (6, 11, 'sp4_r_v_b_10')
// (6, 11, 'sp4_r_v_b_26')
// (6, 11, 'sp4_r_v_b_4')
// (6, 12, 'sp4_r_v_b_15')
// (6, 13, 'sp4_r_v_b_2')
// (7, 7, 'sp4_v_t_41')
// (7, 7, 'sp4_v_t_47')
// (7, 8, 'local_g3_0')
// (7, 8, 'local_g3_1')
// (7, 8, 'lutff_2/in_2')
// (7, 8, 'lutff_3/in_2')
// (7, 8, 'lutff_4/in_0')
// (7, 8, 'sp4_h_r_32')
// (7, 8, 'sp4_v_b_41')
// (7, 8, 'sp4_v_b_47')
// (7, 9, 'sp4_h_l_39')
// (7, 9, 'sp4_v_b_28')
// (7, 9, 'sp4_v_b_34')
// (7, 9, 'sp4_v_t_39')
// (7, 10, 'local_g0_1')
// (7, 10, 'local_g1_7')
// (7, 10, 'lutff_2/in_2')
// (7, 10, 'lutff_3/in_2')
// (7, 10, 'lutff_5/in_2')
// (7, 10, 'lutff_6/in_0')
// (7, 10, 'sp4_v_b_17')
// (7, 10, 'sp4_v_b_23')
// (7, 10, 'sp4_v_b_39')
// (7, 11, 'sp4_h_l_47')
// (7, 11, 'sp4_v_b_10')
// (7, 11, 'sp4_v_b_26')
// (7, 11, 'sp4_v_b_4')
// (7, 12, 'sp4_v_b_15')
// (7, 13, 'sp4_v_b_2')
// (8, 8, 'sp4_h_r_45')
// (9, 8, 'sp4_h_l_45')

wire n63;
// (1, 7, 'sp4_h_r_11')
// (2, 7, 'sp4_h_r_22')
// (3, 7, 'sp4_h_r_35')
// (4, 4, 'sp4_r_v_b_46')
// (4, 5, 'neigh_op_tnr_3')
// (4, 5, 'sp4_r_v_b_35')
// (4, 6, 'local_g2_3')
// (4, 6, 'lutff_1/in_2')
// (4, 6, 'lutff_6/in_1')
// (4, 6, 'neigh_op_rgt_3')
// (4, 6, 'sp4_r_v_b_22')
// (4, 7, 'local_g2_3')
// (4, 7, 'local_g2_6')
// (4, 7, 'lutff_1/in_2')
// (4, 7, 'lutff_2/in_2')
// (4, 7, 'neigh_op_bnr_3')
// (4, 7, 'sp4_h_r_46')
// (4, 7, 'sp4_r_v_b_11')
// (5, 3, 'sp4_v_t_46')
// (5, 4, 'sp4_v_b_46')
// (5, 5, 'neigh_op_top_3')
// (5, 5, 'sp4_v_b_35')
// (5, 6, 'local_g1_3')
// (5, 6, 'lutff_3/out')
// (5, 6, 'lutff_6/in_2')
// (5, 6, 'sp4_v_b_22')
// (5, 7, 'neigh_op_bot_3')
// (5, 7, 'sp4_h_l_46')
// (5, 7, 'sp4_v_b_11')
// (6, 5, 'neigh_op_tnl_3')
// (6, 6, 'neigh_op_lft_3')
// (6, 7, 'neigh_op_bnl_3')

wire n64;
// (1, 8, 'neigh_op_tnr_2')
// (1, 9, 'neigh_op_rgt_2')
// (1, 10, 'neigh_op_bnr_2')
// (2, 6, 'sp4_r_v_b_40')
// (2, 7, 'sp4_r_v_b_29')
// (2, 8, 'neigh_op_top_2')
// (2, 8, 'sp4_r_v_b_16')
// (2, 9, 'lutff_2/out')
// (2, 9, 'sp4_r_v_b_5')
// (2, 10, 'neigh_op_bot_2')
// (3, 5, 'sp4_v_t_40')
// (3, 6, 'sp4_v_b_40')
// (3, 7, 'sp4_v_b_29')
// (3, 8, 'neigh_op_tnl_2')
// (3, 8, 'sp4_v_b_16')
// (3, 9, 'neigh_op_lft_2')
// (3, 9, 'sp4_h_r_11')
// (3, 9, 'sp4_v_b_5')
// (3, 10, 'neigh_op_bnl_2')
// (4, 9, 'sp4_h_r_22')
// (5, 9, 'sp4_h_r_35')
// (6, 9, 'sp4_h_r_46')
// (6, 10, 'sp4_r_v_b_41')
// (6, 11, 'sp4_r_v_b_28')
// (6, 12, 'sp4_r_v_b_17')
// (6, 13, 'sp4_r_v_b_4')
// (7, 9, 'sp4_h_l_46')
// (7, 9, 'sp4_v_t_41')
// (7, 10, 'sp4_v_b_41')
// (7, 11, 'sp4_v_b_28')
// (7, 12, 'local_g0_1')
// (7, 12, 'local_g1_1')
// (7, 12, 'lutff_0/in_1')
// (7, 12, 'lutff_5/in_1')
// (7, 12, 'sp4_v_b_17')
// (7, 13, 'sp4_v_b_4')

reg n65 = 0;
// (1, 8, 'neigh_op_tnr_3')
// (1, 9, 'neigh_op_rgt_3')
// (1, 10, 'neigh_op_bnr_3')
// (2, 8, 'local_g0_3')
// (2, 8, 'lutff_2/in_1')
// (2, 8, 'neigh_op_top_3')
// (2, 9, 'local_g1_3')
// (2, 9, 'lutff_2/in_2')
// (2, 9, 'lutff_3/out')
// (2, 10, 'neigh_op_bot_3')
// (3, 8, 'neigh_op_tnl_3')
// (3, 9, 'neigh_op_lft_3')
// (3, 10, 'neigh_op_bnl_3')

reg n66 = 0;
// (1, 8, 'neigh_op_tnr_4')
// (1, 9, 'neigh_op_rgt_4')
// (1, 10, 'neigh_op_bnr_4')
// (2, 8, 'neigh_op_top_4')
// (2, 9, 'local_g1_4')
// (2, 9, 'lutff_2/in_1')
// (2, 9, 'lutff_4/out')
// (2, 10, 'neigh_op_bot_4')
// (3, 8, 'neigh_op_tnl_4')
// (3, 9, 'neigh_op_lft_4')
// (3, 10, 'neigh_op_bnl_4')

reg n67 = 0;
// (1, 8, 'neigh_op_tnr_7')
// (1, 9, 'neigh_op_rgt_7')
// (1, 10, 'neigh_op_bnr_7')
// (2, 8, 'neigh_op_top_7')
// (2, 9, 'local_g0_7')
// (2, 9, 'lutff_4/in_1')
// (2, 9, 'lutff_7/out')
// (2, 10, 'neigh_op_bot_7')
// (3, 8, 'neigh_op_tnl_7')
// (3, 9, 'neigh_op_lft_7')
// (3, 10, 'neigh_op_bnl_7')

reg n68 = 0;
// (1, 9, 'neigh_op_tnr_2')
// (1, 10, 'neigh_op_rgt_2')
// (1, 10, 'sp4_h_r_9')
// (1, 11, 'neigh_op_bnr_2')
// (2, 9, 'neigh_op_top_2')
// (2, 10, 'lutff_2/out')
// (2, 10, 'sp4_h_r_20')
// (2, 11, 'neigh_op_bot_2')
// (3, 9, 'neigh_op_tnl_2')
// (3, 10, 'neigh_op_lft_2')
// (3, 10, 'sp4_h_r_33')
// (3, 11, 'neigh_op_bnl_2')
// (4, 10, 'local_g2_4')
// (4, 10, 'lutff_7/in_1')
// (4, 10, 'sp4_h_r_44')
// (5, 10, 'sp4_h_l_44')

reg n69 = 0;
// (1, 9, 'neigh_op_tnr_7')
// (1, 10, 'neigh_op_rgt_7')
// (1, 11, 'neigh_op_bnr_7')
// (2, 9, 'local_g1_7')
// (2, 9, 'lutff_7/in_1')
// (2, 9, 'neigh_op_top_7')
// (2, 10, 'lutff_7/out')
// (2, 11, 'neigh_op_bot_7')
// (3, 9, 'neigh_op_tnl_7')
// (3, 10, 'neigh_op_lft_7')
// (3, 11, 'neigh_op_bnl_7')

reg n70 = 0;
// (1, 9, 'sp12_h_r_0')
// (2, 9, 'sp12_h_r_3')
// (3, 9, 'sp12_h_r_4')
// (4, 9, 'sp12_h_r_7')
// (5, 9, 'sp12_h_r_8')
// (6, 9, 'sp12_h_r_11')
// (7, 9, 'sp12_h_r_12')
// (8, 8, 'neigh_op_tnr_4')
// (8, 9, 'neigh_op_rgt_4')
// (8, 9, 'sp12_h_r_15')
// (8, 10, 'neigh_op_bnr_4')
// (9, 8, 'neigh_op_top_4')
// (9, 9, 'lutff_4/out')
// (9, 9, 'sp12_h_r_16')
// (9, 10, 'neigh_op_bot_4')
// (10, 8, 'neigh_op_tnl_4')
// (10, 9, 'neigh_op_lft_4')
// (10, 9, 'sp12_h_r_19')
// (10, 10, 'neigh_op_bnl_4')
// (11, 9, 'local_g0_4')
// (11, 9, 'lutff_4/in_0')
// (11, 9, 'sp12_h_r_20')
// (12, 9, 'sp12_h_r_23')
// (13, 9, 'span12_horz_23')

reg n71 = 0;
// (1, 9, 'sp4_h_r_5')
// (2, 9, 'local_g0_0')
// (2, 9, 'lutff_3/in_1')
// (2, 9, 'lutff_4/in_2')
// (2, 9, 'sp4_h_r_16')
// (3, 8, 'neigh_op_tnr_4')
// (3, 9, 'neigh_op_rgt_4')
// (3, 9, 'sp4_h_r_29')
// (3, 10, 'neigh_op_bnr_4')
// (4, 8, 'neigh_op_top_4')
// (4, 9, 'lutff_4/out')
// (4, 9, 'sp4_h_r_40')
// (4, 10, 'neigh_op_bot_4')
// (5, 8, 'neigh_op_tnl_4')
// (5, 9, 'neigh_op_lft_4')
// (5, 9, 'sp4_h_l_40')
// (5, 10, 'neigh_op_bnl_4')

reg n72 = 0;
// (1, 9, 'sp4_h_r_7')
// (2, 9, 'local_g1_2')
// (2, 9, 'lutff_7/in_2')
// (2, 9, 'sp4_h_r_18')
// (3, 8, 'neigh_op_tnr_5')
// (3, 9, 'neigh_op_rgt_5')
// (3, 9, 'sp4_h_r_31')
// (3, 10, 'neigh_op_bnr_5')
// (4, 8, 'neigh_op_top_5')
// (4, 9, 'local_g0_5')
// (4, 9, 'lutff_4/in_1')
// (4, 9, 'lutff_5/out')
// (4, 9, 'sp4_h_r_42')
// (4, 10, 'neigh_op_bot_5')
// (5, 8, 'neigh_op_tnl_5')
// (5, 9, 'neigh_op_lft_5')
// (5, 9, 'sp4_h_l_42')
// (5, 10, 'neigh_op_bnl_5')

reg n73 = 0;
// (1, 10, 'neigh_op_tnr_0')
// (1, 11, 'neigh_op_rgt_0')
// (1, 12, 'neigh_op_bnr_0')
// (2, 10, 'neigh_op_top_0')
// (2, 11, 'local_g1_0')
// (2, 11, 'lutff_0/out')
// (2, 11, 'lutff_1/in_0')
// (2, 12, 'neigh_op_bot_0')
// (3, 10, 'neigh_op_tnl_0')
// (3, 11, 'neigh_op_lft_0')
// (3, 12, 'neigh_op_bnl_0')

reg n74 = 0;
// (1, 10, 'neigh_op_tnr_1')
// (1, 11, 'neigh_op_rgt_1')
// (1, 12, 'neigh_op_bnr_1')
// (2, 10, 'neigh_op_top_1')
// (2, 11, 'local_g0_1')
// (2, 11, 'lutff_1/out')
// (2, 11, 'lutff_5/in_0')
// (2, 12, 'neigh_op_bot_1')
// (3, 10, 'neigh_op_tnl_1')
// (3, 11, 'neigh_op_lft_1')
// (3, 12, 'neigh_op_bnl_1')

reg n75 = 0;
// (1, 10, 'neigh_op_tnr_3')
// (1, 11, 'neigh_op_rgt_3')
// (1, 12, 'neigh_op_bnr_3')
// (2, 10, 'neigh_op_top_3')
// (2, 11, 'local_g1_3')
// (2, 11, 'lutff_2/in_0')
// (2, 11, 'lutff_3/out')
// (2, 12, 'neigh_op_bot_3')
// (3, 10, 'neigh_op_tnl_3')
// (3, 11, 'neigh_op_lft_3')
// (3, 12, 'neigh_op_bnl_3')

reg n76 = 0;
// (1, 10, 'neigh_op_tnr_5')
// (1, 11, 'neigh_op_rgt_5')
// (1, 11, 'sp12_h_r_1')
// (1, 12, 'neigh_op_bnr_5')
// (2, 10, 'neigh_op_top_5')
// (2, 11, 'lutff_5/out')
// (2, 11, 'sp12_h_r_2')
// (2, 12, 'neigh_op_bot_5')
// (3, 10, 'neigh_op_tnl_5')
// (3, 11, 'neigh_op_lft_5')
// (3, 11, 'sp12_h_r_5')
// (3, 12, 'neigh_op_bnl_5')
// (4, 11, 'sp12_h_r_6')
// (5, 11, 'local_g0_1')
// (5, 11, 'lutff_7/in_0')
// (5, 11, 'sp12_h_r_9')
// (6, 11, 'sp12_h_r_10')
// (7, 11, 'sp12_h_r_13')
// (8, 11, 'sp12_h_r_14')
// (9, 11, 'sp12_h_r_17')
// (10, 11, 'sp12_h_r_18')
// (11, 11, 'sp12_h_r_21')
// (12, 11, 'sp12_h_r_22')
// (13, 11, 'span12_horz_22')

reg n77 = 0;
// (1, 10, 'neigh_op_tnr_6')
// (1, 11, 'neigh_op_rgt_6')
// (1, 12, 'neigh_op_bnr_6')
// (2, 10, 'neigh_op_top_6')
// (2, 11, 'local_g1_6')
// (2, 11, 'lutff_3/in_0')
// (2, 11, 'lutff_6/out')
// (2, 12, 'neigh_op_bot_6')
// (3, 10, 'neigh_op_tnl_6')
// (3, 11, 'neigh_op_lft_6')
// (3, 12, 'neigh_op_bnl_6')

reg n78 = 0;
// (1, 11, 'sp4_h_r_5')
// (2, 11, 'local_g0_0')
// (2, 11, 'lutff_0/in_0')
// (2, 11, 'sp4_h_r_16')
// (3, 11, 'sp4_h_r_29')
// (4, 11, 'sp4_h_r_40')
// (5, 11, 'sp4_h_l_40')
// (5, 11, 'sp4_h_r_2')
// (6, 10, 'neigh_op_tnr_5')
// (6, 11, 'neigh_op_rgt_5')
// (6, 11, 'sp4_h_r_15')
// (6, 12, 'neigh_op_bnr_5')
// (7, 10, 'neigh_op_top_5')
// (7, 11, 'lutff_5/out')
// (7, 11, 'sp4_h_r_26')
// (7, 12, 'neigh_op_bot_5')
// (8, 10, 'neigh_op_tnl_5')
// (8, 11, 'neigh_op_lft_5')
// (8, 11, 'sp4_h_r_39')
// (8, 12, 'neigh_op_bnl_5')
// (9, 11, 'sp4_h_l_39')

reg n79 = 0;
// (1, 12, 'neigh_op_tnr_0')
// (1, 13, 'neigh_op_rgt_0')
// (1, 14, 'neigh_op_bnr_0')
// (2, 12, 'neigh_op_top_0')
// (2, 13, 'local_g1_0')
// (2, 13, 'lutff_0/out')
// (2, 13, 'lutff_7/in_0')
// (2, 14, 'neigh_op_bot_0')
// (3, 12, 'neigh_op_tnl_0')
// (3, 13, 'neigh_op_lft_0')
// (3, 14, 'neigh_op_bnl_0')

reg n80 = 0;
// (1, 12, 'neigh_op_tnr_2')
// (1, 13, 'neigh_op_rgt_2')
// (1, 14, 'neigh_op_bnr_2')
// (2, 12, 'neigh_op_top_2')
// (2, 13, 'local_g1_2')
// (2, 13, 'lutff_2/out')
// (2, 13, 'lutff_5/in_0')
// (2, 14, 'neigh_op_bot_2')
// (3, 12, 'neigh_op_tnl_2')
// (3, 13, 'neigh_op_lft_2')
// (3, 14, 'neigh_op_bnl_2')

reg n81 = 0;
// (1, 12, 'neigh_op_tnr_3')
// (1, 13, 'neigh_op_rgt_3')
// (1, 14, 'neigh_op_bnr_3')
// (2, 12, 'neigh_op_top_3')
// (2, 13, 'local_g1_3')
// (2, 13, 'lutff_3/out')
// (2, 13, 'lutff_4/in_0')
// (2, 14, 'neigh_op_bot_3')
// (3, 12, 'neigh_op_tnl_3')
// (3, 13, 'neigh_op_lft_3')
// (3, 14, 'neigh_op_bnl_3')

reg n82 = 0;
// (1, 12, 'neigh_op_tnr_5')
// (1, 13, 'neigh_op_rgt_5')
// (1, 13, 'sp12_h_r_1')
// (1, 14, 'neigh_op_bnr_5')
// (2, 12, 'neigh_op_top_5')
// (2, 13, 'lutff_5/out')
// (2, 13, 'sp12_h_r_2')
// (2, 14, 'neigh_op_bot_5')
// (3, 12, 'neigh_op_tnl_5')
// (3, 13, 'neigh_op_lft_5')
// (3, 13, 'sp12_h_r_5')
// (3, 14, 'neigh_op_bnl_5')
// (4, 13, 'local_g0_6')
// (4, 13, 'lutff_0/in_0')
// (4, 13, 'lutff_5/in_1')
// (4, 13, 'sp12_h_r_6')
// (5, 13, 'sp12_h_r_9')
// (6, 13, 'sp12_h_r_10')
// (7, 13, 'sp12_h_r_13')
// (8, 13, 'sp12_h_r_14')
// (9, 13, 'sp12_h_r_17')
// (10, 13, 'sp12_h_r_18')
// (11, 13, 'sp12_h_r_21')
// (12, 13, 'sp12_h_r_22')
// (13, 13, 'span12_horz_22')

reg n83 = 0;
// (1, 12, 'neigh_op_tnr_7')
// (1, 13, 'neigh_op_rgt_7')
// (1, 14, 'neigh_op_bnr_7')
// (2, 12, 'neigh_op_top_7')
// (2, 13, 'local_g1_7')
// (2, 13, 'lutff_2/in_0')
// (2, 13, 'lutff_7/out')
// (2, 14, 'neigh_op_bot_7')
// (3, 12, 'neigh_op_tnl_7')
// (3, 13, 'neigh_op_lft_7')
// (3, 14, 'neigh_op_bnl_7')

wire n84;
// (1, 12, 'sp12_h_r_1')
// (2, 12, 'sp12_h_r_2')
// (3, 12, 'sp12_h_r_5')
// (4, 12, 'sp12_h_r_6')
// (5, 11, 'neigh_op_tnr_1')
// (5, 12, 'neigh_op_rgt_1')
// (5, 12, 'sp12_h_r_9')
// (5, 13, 'neigh_op_bnr_1')
// (6, 11, 'neigh_op_top_1')
// (6, 12, 'local_g1_2')
// (6, 12, 'lutff_0/in_3')
// (6, 12, 'lutff_1/out')
// (6, 12, 'sp12_h_r_10')
// (6, 13, 'neigh_op_bot_1')
// (7, 11, 'neigh_op_tnl_1')
// (7, 12, 'neigh_op_lft_1')
// (7, 12, 'sp12_h_r_13')
// (7, 13, 'neigh_op_bnl_1')
// (8, 12, 'sp12_h_r_14')
// (9, 12, 'sp12_h_r_17')
// (10, 12, 'sp12_h_r_18')
// (11, 12, 'sp12_h_r_21')
// (12, 12, 'sp12_h_r_22')
// (13, 12, 'span12_horz_22')

reg n85 = 0;
// (1, 12, 'sp4_h_r_5')
// (2, 12, 'local_g1_0')
// (2, 12, 'lutff_7/in_0')
// (2, 12, 'sp4_h_r_16')
// (3, 11, 'neigh_op_tnr_4')
// (3, 12, 'neigh_op_rgt_4')
// (3, 12, 'sp4_h_r_29')
// (3, 13, 'neigh_op_bnr_4')
// (4, 11, 'neigh_op_top_4')
// (4, 12, 'lutff_4/out')
// (4, 12, 'sp4_h_r_40')
// (4, 13, 'neigh_op_bot_4')
// (5, 11, 'neigh_op_tnl_4')
// (5, 12, 'neigh_op_lft_4')
// (5, 12, 'sp4_h_l_40')
// (5, 13, 'neigh_op_bnl_4')

reg n86 = 0;
// (1, 13, 'neigh_op_tnr_5')
// (1, 14, 'neigh_op_rgt_5')
// (1, 14, 'sp12_h_r_1')
// (1, 15, 'neigh_op_bnr_5')
// (2, 13, 'neigh_op_top_5')
// (2, 14, 'lutff_5/out')
// (2, 14, 'sp12_h_r_2')
// (2, 15, 'neigh_op_bot_5')
// (3, 13, 'neigh_op_tnl_5')
// (3, 14, 'neigh_op_lft_5')
// (3, 14, 'sp12_h_r_5')
// (3, 15, 'neigh_op_bnl_5')
// (4, 14, 'sp12_h_r_6')
// (5, 14, 'local_g0_1')
// (5, 14, 'lutff_5/in_0')
// (5, 14, 'sp12_h_r_9')
// (6, 14, 'sp12_h_r_10')
// (7, 14, 'sp12_h_r_13')
// (8, 14, 'sp12_h_r_14')
// (9, 14, 'sp12_h_r_17')
// (10, 14, 'sp12_h_r_18')
// (11, 14, 'sp12_h_r_21')
// (12, 14, 'sp12_h_r_22')
// (13, 14, 'span12_horz_22')

wire n87;
// (2, 2, 'sp4_h_r_7')
// (3, 2, 'sp4_h_r_18')
// (4, 2, 'sp4_h_r_31')
// (5, 1, 'sp4_r_v_b_18')
// (5, 2, 'sp4_h_r_42')
// (5, 2, 'sp4_r_v_b_7')
// (5, 3, 'sp4_r_v_b_47')
// (5, 4, 'sp4_r_v_b_34')
// (5, 5, 'sp4_r_v_b_23')
// (5, 6, 'sp4_r_v_b_10')
// (6, 0, 'span4_vert_18')
// (6, 1, 'sp4_v_b_18')
// (6, 2, 'local_g1_7')
// (6, 2, 'lutff_3/in_3')
// (6, 2, 'sp4_h_l_42')
// (6, 2, 'sp4_h_r_4')
// (6, 2, 'sp4_v_b_7')
// (6, 2, 'sp4_v_t_47')
// (6, 3, 'local_g2_7')
// (6, 3, 'local_g3_7')
// (6, 3, 'lutff_0/in_1')
// (6, 3, 'lutff_1/in_0')
// (6, 3, 'lutff_2/in_2')
// (6, 3, 'lutff_3/in_3')
// (6, 3, 'lutff_6/in_3')
// (6, 3, 'lutff_7/in_1')
// (6, 3, 'sp4_v_b_47')
// (6, 4, 'sp4_v_b_34')
// (6, 5, 'sp4_v_b_23')
// (6, 6, 'sp4_v_b_10')
// (7, 1, 'neigh_op_tnr_6')
// (7, 2, 'local_g3_6')
// (7, 2, 'lutff_2/in_3')
// (7, 2, 'neigh_op_rgt_6')
// (7, 2, 'sp4_h_r_17')
// (7, 3, 'neigh_op_bnr_6')
// (8, 1, 'neigh_op_top_6')
// (8, 2, 'lutff_6/out')
// (8, 2, 'sp4_h_r_28')
// (8, 3, 'neigh_op_bot_6')
// (9, 1, 'neigh_op_tnl_6')
// (9, 2, 'neigh_op_lft_6')
// (9, 2, 'sp4_h_r_41')
// (9, 3, 'neigh_op_bnl_6')
// (10, 2, 'sp4_h_l_41')

wire n88;
// (2, 3, 'sp12_h_r_0')
// (3, 3, 'sp12_h_r_3')
// (4, 3, 'sp12_h_r_4')
// (5, 2, 'neigh_op_tnr_0')
// (5, 3, 'neigh_op_rgt_0')
// (5, 3, 'sp12_h_r_7')
// (5, 4, 'neigh_op_bnr_0')
// (6, 2, 'neigh_op_top_0')
// (6, 3, 'lutff_0/out')
// (6, 3, 'sp12_h_r_8')
// (6, 4, 'neigh_op_bot_0')
// (7, 2, 'neigh_op_tnl_0')
// (7, 3, 'local_g0_3')
// (7, 3, 'local_g1_3')
// (7, 3, 'lutff_1/in_1')
// (7, 3, 'lutff_6/in_1')
// (7, 3, 'neigh_op_lft_0')
// (7, 3, 'sp12_h_r_11')
// (7, 4, 'neigh_op_bnl_0')
// (8, 3, 'sp12_h_r_12')
// (9, 3, 'sp12_h_r_15')
// (10, 3, 'sp12_h_r_16')
// (11, 3, 'sp12_h_r_19')
// (12, 3, 'sp12_h_r_20')
// (13, 3, 'span12_horz_20')

wire n89;
// (2, 3, 'sp12_h_r_1')
// (3, 3, 'sp12_h_r_2')
// (4, 3, 'sp12_h_r_5')
// (5, 3, 'sp12_h_r_6')
// (6, 3, 'sp12_h_r_9')
// (7, 2, 'local_g0_1')
// (7, 2, 'lutff_1/in_0')
// (7, 2, 'lutff_7/in_0')
// (7, 2, 'sp4_h_r_1')
// (7, 3, 'local_g0_2')
// (7, 3, 'local_g1_2')
// (7, 3, 'lutff_4/in_3')
// (7, 3, 'lutff_7/in_3')
// (7, 3, 'sp12_h_r_10')
// (8, 2, 'local_g0_4')
// (8, 2, 'lutff_6/in_0')
// (8, 2, 'sp4_h_r_12')
// (8, 3, 'sp12_h_r_13')
// (9, 2, 'sp4_h_r_25')
// (9, 3, 'sp12_h_r_14')
// (10, 2, 'neigh_op_tnr_5')
// (10, 2, 'sp4_h_r_36')
// (10, 3, 'neigh_op_rgt_5')
// (10, 3, 'sp12_h_r_17')
// (10, 3, 'sp4_r_v_b_42')
// (10, 4, 'neigh_op_bnr_5')
// (10, 4, 'sp4_r_v_b_31')
// (10, 5, 'sp4_r_v_b_18')
// (10, 6, 'sp4_r_v_b_7')
// (11, 2, 'neigh_op_top_5')
// (11, 2, 'sp4_h_l_36')
// (11, 2, 'sp4_v_t_42')
// (11, 3, 'lutff_5/out')
// (11, 3, 'sp12_h_r_18')
// (11, 3, 'sp4_v_b_42')
// (11, 4, 'neigh_op_bot_5')
// (11, 4, 'sp4_v_b_31')
// (11, 5, 'sp4_v_b_18')
// (11, 6, 'sp4_v_b_7')
// (12, 2, 'neigh_op_tnl_5')
// (12, 3, 'neigh_op_lft_5')
// (12, 3, 'sp12_h_r_21')
// (12, 4, 'neigh_op_bnl_5')
// (13, 3, 'span12_horz_21')

reg n90 = 0;
// (2, 3, 'sp4_r_v_b_39')
// (2, 4, 'local_g0_2')
// (2, 4, 'lutff_4/in_0')
// (2, 4, 'sp4_r_v_b_26')
// (2, 5, 'sp4_r_v_b_15')
// (2, 6, 'sp4_r_v_b_2')
// (3, 2, 'sp4_v_t_39')
// (3, 3, 'sp4_v_b_39')
// (3, 4, 'sp4_v_b_26')
// (3, 5, 'sp4_v_b_15')
// (3, 6, 'sp4_h_r_9')
// (3, 6, 'sp4_v_b_2')
// (3, 12, 'sp4_h_r_4')
// (4, 6, 'sp4_h_r_20')
// (4, 12, 'local_g0_1')
// (4, 12, 'lutff_3/in_0')
// (4, 12, 'sp4_h_r_17')
// (5, 6, 'sp4_h_r_33')
// (5, 12, 'local_g2_4')
// (5, 12, 'local_g3_4')
// (5, 12, 'lutff_0/in_2')
// (5, 12, 'lutff_7/in_2')
// (5, 12, 'sp4_h_r_28')
// (6, 5, 'sp4_r_v_b_46')
// (6, 6, 'neigh_op_tnr_3')
// (6, 6, 'sp4_h_r_44')
// (6, 6, 'sp4_r_v_b_35')
// (6, 7, 'neigh_op_rgt_3')
// (6, 7, 'sp4_r_v_b_22')
// (6, 7, 'sp4_r_v_b_38')
// (6, 8, 'neigh_op_bnr_3')
// (6, 8, 'sp4_r_v_b_11')
// (6, 8, 'sp4_r_v_b_27')
// (6, 9, 'sp4_r_v_b_14')
// (6, 9, 'sp4_r_v_b_46')
// (6, 10, 'sp4_r_v_b_3')
// (6, 10, 'sp4_r_v_b_35')
// (6, 11, 'sp4_r_v_b_22')
// (6, 12, 'sp4_h_r_41')
// (6, 12, 'sp4_r_v_b_11')
// (7, 4, 'sp4_v_t_46')
// (7, 5, 'sp4_v_b_46')
// (7, 6, 'neigh_op_top_3')
// (7, 6, 'sp4_h_l_44')
// (7, 6, 'sp4_v_b_35')
// (7, 6, 'sp4_v_t_38')
// (7, 7, 'lutff_3/out')
// (7, 7, 'sp4_v_b_22')
// (7, 7, 'sp4_v_b_38')
// (7, 8, 'neigh_op_bot_3')
// (7, 8, 'sp4_v_b_11')
// (7, 8, 'sp4_v_b_27')
// (7, 8, 'sp4_v_t_46')
// (7, 9, 'sp4_v_b_14')
// (7, 9, 'sp4_v_b_46')
// (7, 10, 'sp4_v_b_3')
// (7, 10, 'sp4_v_b_35')
// (7, 11, 'sp4_v_b_22')
// (7, 12, 'sp4_h_l_41')
// (7, 12, 'sp4_v_b_11')
// (8, 6, 'neigh_op_tnl_3')
// (8, 7, 'neigh_op_lft_3')
// (8, 8, 'neigh_op_bnl_3')

wire n91;
// (2, 4, 'local_g0_1')
// (2, 4, 'lutff_2/in_1')
// (2, 4, 'sp4_h_r_1')
// (3, 4, 'sp4_h_r_12')
// (4, 3, 'neigh_op_tnr_2')
// (4, 4, 'neigh_op_rgt_2')
// (4, 4, 'sp4_h_r_25')
// (4, 5, 'neigh_op_bnr_2')
// (5, 3, 'neigh_op_top_2')
// (5, 4, 'lutff_2/out')
// (5, 4, 'sp4_h_r_36')
// (5, 5, 'neigh_op_bot_2')
// (6, 3, 'neigh_op_tnl_2')
// (6, 4, 'local_g0_2')
// (6, 4, 'lutff_2/in_2')
// (6, 4, 'lutff_6/in_2')
// (6, 4, 'neigh_op_lft_2')
// (6, 4, 'sp4_h_l_36')
// (6, 5, 'neigh_op_bnl_2')

reg n92 = 0;
// (2, 4, 'sp4_h_r_10')
// (3, 4, 'sp4_h_r_23')
// (4, 1, 'neigh_op_tnr_6')
// (4, 2, 'neigh_op_rgt_6')
// (4, 3, 'neigh_op_bnr_6')
// (4, 4, 'sp4_h_r_34')
// (5, 0, 'span12_vert_15')
// (5, 1, 'neigh_op_top_6')
// (5, 1, 'sp12_v_b_15')
// (5, 1, 'sp4_r_v_b_40')
// (5, 2, 'local_g1_6')
// (5, 2, 'lutff_2/in_3')
// (5, 2, 'lutff_4/in_3')
// (5, 2, 'lutff_6/out')
// (5, 2, 'sp12_v_b_12')
// (5, 2, 'sp4_r_v_b_29')
// (5, 2, 'sp4_r_v_b_45')
// (5, 3, 'neigh_op_bot_6')
// (5, 3, 'sp12_v_b_11')
// (5, 3, 'sp4_r_v_b_16')
// (5, 3, 'sp4_r_v_b_32')
// (5, 4, 'local_g3_0')
// (5, 4, 'lutff_1/in_0')
// (5, 4, 'sp12_v_b_8')
// (5, 4, 'sp4_h_r_47')
// (5, 4, 'sp4_r_v_b_21')
// (5, 4, 'sp4_r_v_b_5')
// (5, 5, 'sp12_v_b_7')
// (5, 5, 'sp4_r_v_b_8')
// (5, 6, 'sp12_v_b_4')
// (5, 7, 'sp12_v_b_3')
// (5, 8, 'sp12_v_b_0')
// (6, 0, 'span4_vert_40')
// (6, 1, 'neigh_op_tnl_6')
// (6, 1, 'sp4_v_b_40')
// (6, 1, 'sp4_v_t_45')
// (6, 2, 'neigh_op_lft_6')
// (6, 2, 'sp4_v_b_29')
// (6, 2, 'sp4_v_b_45')
// (6, 3, 'neigh_op_bnl_6')
// (6, 3, 'sp4_v_b_16')
// (6, 3, 'sp4_v_b_32')
// (6, 4, 'local_g0_3')
// (6, 4, 'lutff_3/in_2')
// (6, 4, 'sp4_h_l_47')
// (6, 4, 'sp4_h_r_1')
// (6, 4, 'sp4_h_r_11')
// (6, 4, 'sp4_v_b_21')
// (6, 4, 'sp4_v_b_5')
// (6, 5, 'sp4_h_r_1')
// (6, 5, 'sp4_h_r_2')
// (6, 5, 'sp4_v_b_8')
// (6, 8, 'sp4_h_r_9')
// (7, 4, 'local_g1_4')
// (7, 4, 'lutff_7/in_0')
// (7, 4, 'sp4_h_r_12')
// (7, 4, 'sp4_h_r_22')
// (7, 5, 'local_g1_7')
// (7, 5, 'lutff_4/in_0')
// (7, 5, 'sp4_h_r_12')
// (7, 5, 'sp4_h_r_15')
// (7, 8, 'sp4_h_r_20')
// (8, 4, 'sp4_h_r_25')
// (8, 4, 'sp4_h_r_35')
// (8, 5, 'local_g2_1')
// (8, 5, 'local_g2_2')
// (8, 5, 'lutff_1/in_0')
// (8, 5, 'lutff_4/in_0')
// (8, 5, 'lutff_6/in_0')
// (8, 5, 'sp4_h_r_25')
// (8, 5, 'sp4_h_r_26')
// (8, 8, 'sp4_h_r_33')
// (9, 4, 'local_g3_6')
// (9, 4, 'lutff_5/in_0')
// (9, 4, 'sp4_h_r_36')
// (9, 4, 'sp4_h_r_46')
// (9, 5, 'local_g3_1')
// (9, 5, 'local_g3_4')
// (9, 5, 'lutff_1/in_1')
// (9, 5, 'lutff_4/in_0')
// (9, 5, 'lutff_5/in_0')
// (9, 5, 'sp4_h_r_36')
// (9, 5, 'sp4_h_r_39')
// (9, 5, 'sp4_r_v_b_41')
// (9, 5, 'sp4_r_v_b_44')
// (9, 6, 'sp4_r_v_b_28')
// (9, 6, 'sp4_r_v_b_33')
// (9, 7, 'sp4_r_v_b_17')
// (9, 7, 'sp4_r_v_b_20')
// (9, 8, 'local_g2_4')
// (9, 8, 'lutff_0/in_2')
// (9, 8, 'sp4_h_r_44')
// (9, 8, 'sp4_r_v_b_4')
// (9, 8, 'sp4_r_v_b_9')
// (10, 4, 'sp4_h_l_36')
// (10, 4, 'sp4_h_l_46')
// (10, 4, 'sp4_h_r_7')
// (10, 4, 'sp4_v_t_41')
// (10, 4, 'sp4_v_t_44')
// (10, 5, 'sp4_h_l_36')
// (10, 5, 'sp4_h_l_39')
// (10, 5, 'sp4_h_r_5')
// (10, 5, 'sp4_v_b_41')
// (10, 5, 'sp4_v_b_44')
// (10, 6, 'sp4_v_b_28')
// (10, 6, 'sp4_v_b_33')
// (10, 7, 'sp4_v_b_17')
// (10, 7, 'sp4_v_b_20')
// (10, 8, 'sp4_h_l_44')
// (10, 8, 'sp4_v_b_4')
// (10, 8, 'sp4_v_b_9')
// (11, 4, 'local_g0_2')
// (11, 4, 'lutff_2/in_0')
// (11, 4, 'lutff_6/in_0')
// (11, 4, 'sp4_h_r_18')
// (11, 5, 'local_g0_0')
// (11, 5, 'local_g1_0')
// (11, 5, 'lutff_0/in_0')
// (11, 5, 'lutff_1/in_0')
// (11, 5, 'lutff_3/in_0')
// (11, 5, 'sp4_h_r_16')
// (12, 4, 'sp4_h_r_31')
// (12, 5, 'sp4_h_r_29')
// (13, 4, 'span4_horz_31')
// (13, 5, 'span4_horz_29')

wire n93;
// (2, 5, 'lutff_1/cout')
// (2, 5, 'lutff_2/in_3')

wire n94;
// (2, 5, 'lutff_2/cout')
// (2, 5, 'lutff_3/in_3')

wire n95;
// (2, 5, 'lutff_3/cout')
// (2, 5, 'lutff_4/in_3')

wire n96;
// (2, 5, 'lutff_4/cout')
// (2, 5, 'lutff_5/in_3')

wire n97;
// (2, 5, 'lutff_5/cout')
// (2, 5, 'lutff_6/in_3')

wire n98;
// (2, 5, 'lutff_6/cout')
// (2, 5, 'lutff_7/in_3')

reg n99 = 0;
// (2, 5, 'sp12_h_r_1')
// (3, 5, 'sp12_h_r_2')
// (4, 5, 'sp12_h_r_5')
// (5, 5, 'sp12_h_r_6')
// (6, 5, 'sp12_h_r_9')
// (6, 5, 'sp4_h_r_4')
// (7, 5, 'local_g0_1')
// (7, 5, 'lutff_7/in_0')
// (7, 5, 'sp12_h_r_10')
// (7, 5, 'sp4_h_r_17')
// (8, 5, 'sp12_h_r_13')
// (8, 5, 'sp4_h_r_28')
// (9, 5, 'sp12_h_r_14')
// (9, 5, 'sp4_h_r_41')
// (10, 4, 'neigh_op_tnr_5')
// (10, 5, 'neigh_op_rgt_5')
// (10, 5, 'sp12_h_r_17')
// (10, 5, 'sp4_h_l_41')
// (10, 6, 'neigh_op_bnr_5')
// (11, 4, 'neigh_op_top_5')
// (11, 5, 'lutff_5/out')
// (11, 5, 'sp12_h_r_18')
// (11, 6, 'neigh_op_bot_5')
// (12, 4, 'neigh_op_tnl_5')
// (12, 5, 'neigh_op_lft_5')
// (12, 5, 'sp12_h_r_21')
// (12, 6, 'neigh_op_bnl_5')
// (13, 5, 'span12_horz_21')

wire select;
// (2, 5, 'sp4_h_r_1')
// (3, 5, 'sp4_h_r_12')
// (4, 5, 'local_g2_1')
// (4, 5, 'lutff_4/in_3')
// (4, 5, 'sp4_h_r_25')
// (5, 4, 'sp4_r_v_b_36')
// (5, 4, 'sp4_r_v_b_45')
// (5, 5, 'local_g0_3')
// (5, 5, 'lutff_2/in_3')
// (5, 5, 'sp4_h_r_36')
// (5, 5, 'sp4_r_v_b_25')
// (5, 5, 'sp4_r_v_b_32')
// (5, 6, 'sp4_r_v_b_12')
// (5, 6, 'sp4_r_v_b_21')
// (5, 7, 'sp4_r_v_b_1')
// (5, 7, 'sp4_r_v_b_8')
// (6, 3, 'sp4_v_t_36')
// (6, 3, 'sp4_v_t_45')
// (6, 4, 'sp4_v_b_36')
// (6, 4, 'sp4_v_b_45')
// (6, 5, 'sp4_h_l_36')
// (6, 5, 'sp4_h_r_10')
// (6, 5, 'sp4_v_b_25')
// (6, 5, 'sp4_v_b_32')
// (6, 6, 'local_g0_4')
// (6, 6, 'lutff_3/in_3')
// (6, 6, 'sp4_v_b_12')
// (6, 6, 'sp4_v_b_21')
// (6, 7, 'sp4_h_r_8')
// (6, 7, 'sp4_v_b_1')
// (6, 7, 'sp4_v_b_8')
// (7, 5, 'sp4_h_r_23')
// (7, 7, 'sp4_h_r_21')
// (8, 5, 'sp4_h_r_34')
// (8, 7, 'sp4_h_r_32')
// (9, 5, 'sp4_h_r_47')
// (9, 6, 'sp4_r_v_b_47')
// (9, 7, 'sp4_h_r_45')
// (9, 7, 'sp4_r_v_b_34')
// (9, 8, 'local_g3_5')
// (9, 8, 'lutff_1/in_3')
// (9, 8, 'sp4_r_v_b_23')
// (9, 8, 'sp4_r_v_b_45')
// (9, 9, 'sp4_r_v_b_10')
// (9, 9, 'sp4_r_v_b_32')
// (9, 10, 'sp4_r_v_b_21')
// (9, 11, 'sp4_r_v_b_8')
// (9, 16, 'neigh_op_tnr_2')
// (9, 16, 'neigh_op_tnr_6')
// (10, 5, 'sp4_h_l_47')
// (10, 5, 'sp4_v_t_47')
// (10, 6, 'sp4_v_b_47')
// (10, 7, 'sp12_h_r_0')
// (10, 7, 'sp12_v_t_23')
// (10, 7, 'sp4_h_l_45')
// (10, 7, 'sp4_v_b_34')
// (10, 7, 'sp4_v_t_45')
// (10, 8, 'sp12_v_b_23')
// (10, 8, 'sp4_r_v_b_44')
// (10, 8, 'sp4_v_b_23')
// (10, 8, 'sp4_v_b_45')
// (10, 9, 'sp12_v_b_20')
// (10, 9, 'sp4_h_r_4')
// (10, 9, 'sp4_r_v_b_33')
// (10, 9, 'sp4_v_b_10')
// (10, 9, 'sp4_v_b_32')
// (10, 10, 'sp12_v_b_19')
// (10, 10, 'sp4_r_v_b_20')
// (10, 10, 'sp4_v_b_21')
// (10, 11, 'sp12_v_b_16')
// (10, 11, 'sp4_h_r_8')
// (10, 11, 'sp4_r_v_b_9')
// (10, 11, 'sp4_v_b_8')
// (10, 12, 'sp12_v_b_15')
// (10, 13, 'sp12_v_b_12')
// (10, 14, 'sp12_v_b_11')
// (10, 15, 'sp12_v_b_8')
// (10, 16, 'neigh_op_top_2')
// (10, 16, 'neigh_op_top_6')
// (10, 16, 'sp12_v_b_7')
// (10, 17, 'io_1/D_IN_0')
// (10, 17, 'io_1/PAD')
// (10, 17, 'span12_vert_4')
// (11, 7, 'sp12_h_r_3')
// (11, 7, 'sp4_h_r_3')
// (11, 7, 'sp4_v_t_44')
// (11, 8, 'sp4_v_b_44')
// (11, 9, 'local_g1_1')
// (11, 9, 'lutff_1/in_3')
// (11, 9, 'sp4_h_r_17')
// (11, 9, 'sp4_v_b_33')
// (11, 10, 'local_g0_4')
// (11, 10, 'lutff_1/in_3')
// (11, 10, 'sp4_v_b_20')
// (11, 11, 'local_g1_5')
// (11, 11, 'lutff_1/in_3')
// (11, 11, 'lutff_3/in_3')
// (11, 11, 'sp4_h_r_21')
// (11, 11, 'sp4_v_b_9')
// (11, 16, 'neigh_op_tnl_2')
// (11, 16, 'neigh_op_tnl_6')
// (12, 7, 'sp12_h_r_4')
// (12, 7, 'sp4_h_r_14')
// (12, 9, 'sp4_h_r_28')
// (12, 11, 'sp4_h_r_32')
// (13, 7, 'span12_horz_4')
// (13, 7, 'span4_horz_14')
// (13, 9, 'span4_horz_28')
// (13, 11, 'span4_horz_32')

wire n101;
// (2, 6, 'local_g1_1')
// (2, 6, 'lutff_3/in_3')
// (2, 6, 'sp4_h_r_9')
// (3, 6, 'sp4_h_r_20')
// (4, 5, 'neigh_op_tnr_6')
// (4, 6, 'neigh_op_rgt_6')
// (4, 6, 'sp4_h_r_33')
// (4, 7, 'neigh_op_bnr_6')
// (5, 5, 'neigh_op_top_6')
// (5, 6, 'lutff_6/out')
// (5, 6, 'sp4_h_r_44')
// (5, 7, 'neigh_op_bot_6')
// (6, 5, 'neigh_op_tnl_6')
// (6, 6, 'neigh_op_lft_6')
// (6, 6, 'sp4_h_l_44')
// (6, 7, 'neigh_op_bnl_6')

reg n102 = 0;
// (2, 6, 'sp12_h_r_0')
// (3, 6, 'sp12_h_r_3')
// (4, 6, 'sp12_h_r_4')
// (4, 10, 'sp4_r_v_b_40')
// (4, 11, 'sp4_h_r_10')
// (4, 11, 'sp4_r_v_b_29')
// (4, 12, 'sp4_r_v_b_16')
// (4, 13, 'sp4_r_v_b_5')
// (5, 6, 'sp12_h_r_7')
// (5, 9, 'sp4_h_r_5')
// (5, 9, 'sp4_v_t_40')
// (5, 10, 'sp4_v_b_40')
// (5, 11, 'local_g1_7')
// (5, 11, 'lutff_2/in_2')
// (5, 11, 'sp4_h_r_23')
// (5, 11, 'sp4_v_b_29')
// (5, 12, 'local_g0_0')
// (5, 12, 'lutff_6/in_2')
// (5, 12, 'sp4_v_b_16')
// (5, 13, 'sp4_v_b_5')
// (6, 6, 'sp12_h_r_8')
// (6, 9, 'sp4_h_r_16')
// (6, 11, 'sp4_h_r_34')
// (7, 4, 'sp4_r_v_b_44')
// (7, 5, 'neigh_op_tnr_2')
// (7, 5, 'sp4_r_v_b_33')
// (7, 6, 'neigh_op_rgt_2')
// (7, 6, 'sp12_h_r_11')
// (7, 6, 'sp4_h_r_7')
// (7, 6, 'sp4_r_v_b_20')
// (7, 7, 'neigh_op_bnr_2')
// (7, 7, 'sp4_r_v_b_9')
// (7, 8, 'sp4_r_v_b_40')
// (7, 9, 'sp4_h_r_29')
// (7, 9, 'sp4_r_v_b_29')
// (7, 10, 'sp4_r_v_b_16')
// (7, 11, 'sp4_h_r_47')
// (7, 11, 'sp4_r_v_b_5')
// (8, 3, 'sp4_v_t_44')
// (8, 4, 'sp4_v_b_44')
// (8, 5, 'neigh_op_top_2')
// (8, 5, 'sp4_v_b_33')
// (8, 6, 'lutff_2/out')
// (8, 6, 'sp12_h_r_12')
// (8, 6, 'sp4_h_r_18')
// (8, 6, 'sp4_r_v_b_37')
// (8, 6, 'sp4_v_b_20')
// (8, 7, 'neigh_op_bot_2')
// (8, 7, 'sp4_r_v_b_24')
// (8, 7, 'sp4_v_b_9')
// (8, 7, 'sp4_v_t_40')
// (8, 8, 'sp4_r_v_b_13')
// (8, 8, 'sp4_v_b_40')
// (8, 9, 'sp4_h_r_40')
// (8, 9, 'sp4_r_v_b_0')
// (8, 9, 'sp4_v_b_29')
// (8, 10, 'sp4_v_b_16')
// (8, 11, 'sp4_h_l_47')
// (8, 11, 'sp4_v_b_5')
// (9, 5, 'neigh_op_tnl_2')
// (9, 5, 'sp4_v_t_37')
// (9, 6, 'neigh_op_lft_2')
// (9, 6, 'sp12_h_r_15')
// (9, 6, 'sp4_h_r_31')
// (9, 6, 'sp4_v_b_37')
// (9, 7, 'neigh_op_bnl_2')
// (9, 7, 'sp4_v_b_24')
// (9, 8, 'sp4_v_b_13')
// (9, 9, 'sp4_h_l_40')
// (9, 9, 'sp4_v_b_0')
// (10, 6, 'sp12_h_r_16')
// (10, 6, 'sp4_h_r_42')
// (10, 7, 'sp4_r_v_b_37')
// (10, 8, 'sp4_r_v_b_24')
// (10, 9, 'sp4_r_v_b_13')
// (10, 10, 'sp4_r_v_b_0')
// (11, 6, 'local_g1_3')
// (11, 6, 'lutff_6/in_0')
// (11, 6, 'sp12_h_r_19')
// (11, 6, 'sp4_h_l_42')
// (11, 6, 'sp4_v_t_37')
// (11, 7, 'local_g2_5')
// (11, 7, 'lutff_3/in_0')
// (11, 7, 'sp4_v_b_37')
// (11, 8, 'sp4_v_b_24')
// (11, 9, 'sp4_v_b_13')
// (11, 10, 'sp4_v_b_0')
// (12, 6, 'sp12_h_r_20')
// (13, 6, 'span12_horz_20')

wire n103;
// (2, 7, 'sp4_h_r_3')
// (3, 7, 'sp4_h_r_14')
// (4, 7, 'sp4_h_r_27')
// (5, 7, 'local_g3_6')
// (5, 7, 'lutff_0/in_3')
// (5, 7, 'sp4_h_r_38')
// (5, 8, 'sp4_r_v_b_38')
// (5, 9, 'local_g0_3')
// (5, 9, 'lutff_4/in_3')
// (5, 9, 'sp4_r_v_b_27')
// (5, 10, 'neigh_op_tnr_1')
// (5, 10, 'sp4_r_v_b_14')
// (5, 11, 'neigh_op_rgt_1')
// (5, 11, 'sp4_r_v_b_3')
// (5, 12, 'neigh_op_bnr_1')
// (6, 0, 'span12_vert_22')
// (6, 1, 'sp12_v_b_22')
// (6, 2, 'sp12_v_b_21')
// (6, 3, 'sp12_v_b_18')
// (6, 4, 'sp12_v_b_17')
// (6, 5, 'sp12_v_b_14')
// (6, 6, 'sp12_v_b_13')
// (6, 7, 'local_g3_2')
// (6, 7, 'lutff_2/in_3')
// (6, 7, 'sp12_v_b_10')
// (6, 7, 'sp4_h_l_38')
// (6, 7, 'sp4_v_t_38')
// (6, 8, 'sp12_v_b_9')
// (6, 8, 'sp4_v_b_38')
// (6, 9, 'sp12_v_b_6')
// (6, 9, 'sp4_v_b_27')
// (6, 10, 'neigh_op_top_1')
// (6, 10, 'sp12_v_b_5')
// (6, 10, 'sp4_v_b_14')
// (6, 11, 'lutff_1/out')
// (6, 11, 'sp12_v_b_2')
// (6, 11, 'sp4_v_b_3')
// (6, 12, 'neigh_op_bot_1')
// (6, 12, 'sp12_v_b_1')
// (7, 10, 'neigh_op_tnl_1')
// (7, 11, 'neigh_op_lft_1')
// (7, 12, 'neigh_op_bnl_1')

wire n104;
// (2, 8, 'sp4_h_r_2')
// (3, 7, 'neigh_op_tnr_5')
// (3, 7, 'sp4_r_v_b_39')
// (3, 8, 'neigh_op_rgt_5')
// (3, 8, 'sp4_h_r_15')
// (3, 8, 'sp4_r_v_b_26')
// (3, 8, 'sp4_r_v_b_42')
// (3, 9, 'neigh_op_bnr_5')
// (3, 9, 'sp4_r_v_b_15')
// (3, 9, 'sp4_r_v_b_31')
// (3, 10, 'sp4_r_v_b_18')
// (3, 10, 'sp4_r_v_b_2')
// (3, 11, 'sp4_r_v_b_7')
// (4, 5, 'sp4_r_v_b_46')
// (4, 6, 'sp4_r_v_b_35')
// (4, 6, 'sp4_v_t_39')
// (4, 7, 'neigh_op_top_5')
// (4, 7, 'sp4_r_v_b_22')
// (4, 7, 'sp4_v_b_39')
// (4, 7, 'sp4_v_t_42')
// (4, 8, 'lutff_5/out')
// (4, 8, 'sp4_h_r_26')
// (4, 8, 'sp4_r_v_b_11')
// (4, 8, 'sp4_v_b_26')
// (4, 8, 'sp4_v_b_42')
// (4, 9, 'local_g1_5')
// (4, 9, 'lutff_1/in_3')
// (4, 9, 'neigh_op_bot_5')
// (4, 9, 'sp4_v_b_15')
// (4, 9, 'sp4_v_b_31')
// (4, 10, 'local_g1_2')
// (4, 10, 'lutff_0/in_3')
// (4, 10, 'sp4_v_b_18')
// (4, 10, 'sp4_v_b_2')
// (4, 11, 'local_g1_7')
// (4, 11, 'lutff_3/in_3')
// (4, 11, 'lutff_5/in_3')
// (4, 11, 'sp4_v_b_7')
// (5, 4, 'sp4_v_t_46')
// (5, 5, 'local_g2_6')
// (5, 5, 'lutff_7/in_3')
// (5, 5, 'sp4_v_b_46')
// (5, 6, 'sp4_v_b_35')
// (5, 7, 'neigh_op_tnl_5')
// (5, 7, 'sp4_v_b_22')
// (5, 8, 'neigh_op_lft_5')
// (5, 8, 'sp4_h_r_39')
// (5, 8, 'sp4_v_b_11')
// (5, 9, 'neigh_op_bnl_5')
// (5, 9, 'sp4_r_v_b_42')
// (5, 10, 'sp4_r_v_b_31')
// (5, 11, 'sp4_r_v_b_18')
// (5, 12, 'sp4_r_v_b_7')
// (6, 8, 'sp4_h_l_39')
// (6, 8, 'sp4_v_t_42')
// (6, 9, 'local_g2_2')
// (6, 9, 'lutff_5/in_3')
// (6, 9, 'sp4_v_b_42')
// (6, 10, 'sp4_v_b_31')
// (6, 11, 'sp4_v_b_18')
// (6, 12, 'sp4_v_b_7')

wire n105;
// (2, 9, 'local_g0_2')
// (2, 9, 'lutff_3/in_3')
// (2, 9, 'sp4_h_r_10')
// (3, 8, 'neigh_op_tnr_1')
// (3, 9, 'neigh_op_rgt_1')
// (3, 9, 'sp4_h_r_23')
// (3, 10, 'neigh_op_bnr_1')
// (4, 8, 'neigh_op_top_1')
// (4, 9, 'local_g2_1')
// (4, 9, 'lutff_1/out')
// (4, 9, 'lutff_2/in_3')
// (4, 9, 'lutff_4/in_3')
// (4, 9, 'sp4_h_r_34')
// (4, 10, 'neigh_op_bot_1')
// (5, 6, 'sp4_r_v_b_47')
// (5, 7, 'sp4_r_v_b_34')
// (5, 8, 'neigh_op_tnl_1')
// (5, 8, 'sp4_r_v_b_23')
// (5, 9, 'neigh_op_lft_1')
// (5, 9, 'sp4_h_r_47')
// (5, 9, 'sp4_r_v_b_10')
// (5, 10, 'neigh_op_bnl_1')
// (6, 5, 'sp4_v_t_47')
// (6, 6, 'sp4_v_b_47')
// (6, 7, 'sp4_v_b_34')
// (6, 8, 'sp4_v_b_23')
// (6, 9, 'local_g0_2')
// (6, 9, 'lutff_2/in_2')
// (6, 9, 'sp4_h_l_47')
// (6, 9, 'sp4_h_r_10')
// (6, 9, 'sp4_v_b_10')
// (7, 9, 'sp4_h_r_23')
// (8, 9, 'sp4_h_r_34')
// (9, 9, 'sp4_h_r_47')
// (10, 9, 'sp4_h_l_47')
// (10, 9, 'sp4_h_r_6')
// (11, 9, 'local_g0_3')
// (11, 9, 'lutff_6/in_3')
// (11, 9, 'sp4_h_r_19')
// (12, 9, 'sp4_h_r_30')
// (13, 9, 'span4_horz_30')

reg n106 = 0;
// (2, 9, 'sp12_h_r_1')
// (3, 9, 'sp12_h_r_2')
// (4, 8, 'neigh_op_tnr_7')
// (4, 9, 'neigh_op_rgt_7')
// (4, 9, 'sp12_h_r_5')
// (4, 10, 'neigh_op_bnr_7')
// (5, 8, 'neigh_op_top_7')
// (5, 9, 'lutff_7/out')
// (5, 9, 'sp12_h_r_6')
// (5, 10, 'neigh_op_bot_7')
// (6, 8, 'neigh_op_tnl_7')
// (6, 9, 'local_g0_1')
// (6, 9, 'lutff_6/in_1')
// (6, 9, 'neigh_op_lft_7')
// (6, 9, 'sp12_h_r_9')
// (6, 10, 'neigh_op_bnl_7')
// (7, 9, 'sp12_h_r_10')
// (8, 9, 'sp12_h_r_13')
// (9, 9, 'sp12_h_r_14')
// (10, 9, 'sp12_h_r_17')
// (11, 9, 'sp12_h_r_18')
// (12, 9, 'sp12_h_r_21')
// (13, 9, 'span12_horz_21')

wire n107;
// (2, 9, 'sp4_h_r_11')
// (3, 9, 'sp4_h_r_22')
// (4, 6, 'sp4_h_r_10')
// (4, 6, 'sp4_h_r_4')
// (4, 9, 'sp4_h_r_35')
// (5, 6, 'local_g0_7')
// (5, 6, 'local_g1_1')
// (5, 6, 'lutff_0/in_3')
// (5, 6, 'lutff_7/in_3')
// (5, 6, 'sp4_h_r_17')
// (5, 6, 'sp4_h_r_23')
// (5, 6, 'sp4_r_v_b_40')
// (5, 7, 'local_g0_5')
// (5, 7, 'lutff_2/in_1')
// (5, 7, 'lutff_5/in_2')
// (5, 7, 'sp4_r_v_b_29')
// (5, 8, 'sp4_r_v_b_16')
// (5, 9, 'sp4_h_r_46')
// (5, 9, 'sp4_r_v_b_5')
// (6, 5, 'sp4_v_t_40')
// (6, 6, 'sp4_h_r_28')
// (6, 6, 'sp4_h_r_34')
// (6, 6, 'sp4_v_b_40')
// (6, 7, 'sp4_v_b_29')
// (6, 8, 'neigh_op_tnr_3')
// (6, 8, 'sp4_v_b_16')
// (6, 9, 'neigh_op_rgt_3')
// (6, 9, 'sp4_h_l_46')
// (6, 9, 'sp4_h_r_11')
// (6, 9, 'sp4_v_b_5')
// (6, 10, 'neigh_op_bnr_3')
// (7, 6, 'sp4_h_r_41')
// (7, 6, 'sp4_h_r_47')
// (7, 7, 'sp4_r_v_b_47')
// (7, 8, 'neigh_op_top_3')
// (7, 8, 'sp4_r_v_b_34')
// (7, 9, 'lutff_3/out')
// (7, 9, 'sp4_h_r_22')
// (7, 9, 'sp4_r_v_b_23')
// (7, 10, 'neigh_op_bot_3')
// (7, 10, 'sp4_r_v_b_10')
// (8, 6, 'sp4_h_l_41')
// (8, 6, 'sp4_h_l_47')
// (8, 6, 'sp4_v_t_47')
// (8, 7, 'sp4_v_b_47')
// (8, 8, 'neigh_op_tnl_3')
// (8, 8, 'sp4_v_b_34')
// (8, 9, 'neigh_op_lft_3')
// (8, 9, 'sp4_h_r_35')
// (8, 9, 'sp4_v_b_23')
// (8, 10, 'neigh_op_bnl_3')
// (8, 10, 'sp4_v_b_10')
// (9, 9, 'sp4_h_r_46')
// (10, 9, 'sp4_h_l_46')

reg n108 = 0;
// (2, 11, 'local_g1_1')
// (2, 11, 'lutff_6/in_0')
// (2, 11, 'sp4_h_r_9')
// (3, 11, 'sp4_h_r_20')
// (4, 10, 'neigh_op_tnr_6')
// (4, 11, 'neigh_op_rgt_6')
// (4, 11, 'sp4_h_r_33')
// (4, 12, 'neigh_op_bnr_6')
// (5, 10, 'neigh_op_top_6')
// (5, 11, 'lutff_6/out')
// (5, 11, 'sp4_h_r_44')
// (5, 12, 'neigh_op_bot_6')
// (6, 10, 'neigh_op_tnl_6')
// (6, 11, 'neigh_op_lft_6')
// (6, 11, 'sp4_h_l_44')
// (6, 12, 'neigh_op_bnl_6')

reg n109 = 0;
// (2, 12, 'sp12_h_r_1')
// (3, 12, 'sp12_h_r_2')
// (4, 12, 'sp12_h_r_5')
// (5, 12, 'sp12_h_r_6')
// (6, 11, 'neigh_op_tnr_1')
// (6, 12, 'local_g0_1')
// (6, 12, 'lutff_1/in_0')
// (6, 12, 'neigh_op_rgt_1')
// (6, 12, 'sp12_h_r_9')
// (6, 13, 'local_g0_1')
// (6, 13, 'lutff_2/in_1')
// (6, 13, 'neigh_op_bnr_1')
// (7, 11, 'neigh_op_top_1')
// (7, 12, 'lutff_1/out')
// (7, 12, 'sp12_h_r_10')
// (7, 13, 'neigh_op_bot_1')
// (8, 11, 'neigh_op_tnl_1')
// (8, 12, 'neigh_op_lft_1')
// (8, 12, 'sp12_h_r_13')
// (8, 13, 'neigh_op_bnl_1')
// (9, 12, 'sp12_h_r_14')
// (10, 12, 'sp12_h_r_17')
// (11, 12, 'sp12_h_r_18')
// (12, 12, 'sp12_h_r_21')
// (13, 12, 'span12_horz_21')

reg n110 = 0;
// (2, 13, 'sp12_h_r_1')
// (3, 13, 'sp12_h_r_2')
// (4, 13, 'sp12_h_r_5')
// (5, 13, 'sp12_h_r_6')
// (6, 13, 'sp12_h_r_9')
// (6, 13, 'sp4_h_r_4')
// (7, 13, 'local_g0_1')
// (7, 13, 'lutff_4/in_1')
// (7, 13, 'sp12_h_r_10')
// (7, 13, 'sp4_h_r_17')
// (8, 13, 'local_g2_4')
// (8, 13, 'lutff_1/in_1')
// (8, 13, 'sp12_h_r_13')
// (8, 13, 'sp4_h_r_28')
// (9, 13, 'sp12_h_r_14')
// (9, 13, 'sp4_h_r_41')
// (10, 12, 'neigh_op_tnr_5')
// (10, 13, 'neigh_op_rgt_5')
// (10, 13, 'sp12_h_r_17')
// (10, 13, 'sp4_h_l_41')
// (10, 14, 'neigh_op_bnr_5')
// (11, 12, 'neigh_op_top_5')
// (11, 13, 'lutff_5/out')
// (11, 13, 'sp12_h_r_18')
// (11, 14, 'neigh_op_bot_5')
// (12, 12, 'neigh_op_tnl_5')
// (12, 13, 'neigh_op_lft_5')
// (12, 13, 'sp12_h_r_21')
// (12, 14, 'neigh_op_bnl_5')
// (13, 13, 'span12_horz_21')

reg n111 = 0;
// (2, 14, 'sp12_h_r_0')
// (3, 13, 'neigh_op_tnr_6')
// (3, 14, 'neigh_op_rgt_6')
// (3, 14, 'sp12_h_r_3')
// (3, 15, 'neigh_op_bnr_6')
// (4, 13, 'neigh_op_top_6')
// (4, 14, 'lutff_6/out')
// (4, 14, 'sp12_h_r_4')
// (4, 15, 'neigh_op_bot_6')
// (5, 13, 'neigh_op_tnl_6')
// (5, 14, 'neigh_op_lft_6')
// (5, 14, 'sp12_h_r_7')
// (5, 15, 'neigh_op_bnl_6')
// (6, 14, 'local_g0_0')
// (6, 14, 'local_g1_0')
// (6, 14, 'lutff_0/in_1')
// (6, 14, 'lutff_3/in_1')
// (6, 14, 'sp12_h_r_8')
// (7, 14, 'sp12_h_r_11')
// (8, 14, 'sp12_h_r_12')
// (9, 14, 'sp12_h_r_15')
// (10, 14, 'sp12_h_r_16')
// (11, 14, 'sp12_h_r_19')
// (12, 14, 'sp12_h_r_20')
// (13, 14, 'span12_horz_20')

wire \d_out[5] ;
// (3, 0, 'span4_horz_r_0')
// (4, 0, 'span4_horz_r_4')
// (5, 0, 'io_0/D_OUT_0')
// (5, 0, 'io_0/PAD')
// (5, 0, 'local_g0_0')
// (5, 0, 'span4_horz_r_8')
// (5, 5, 'neigh_op_tnr_3')
// (5, 6, 'neigh_op_rgt_3')
// (5, 7, 'neigh_op_bnr_3')
// (6, 0, 'span4_horz_r_12')
// (6, 1, 'sp4_r_v_b_25')
// (6, 2, 'sp4_r_v_b_12')
// (6, 3, 'sp4_r_v_b_1')
// (6, 4, 'sp4_r_v_b_47')
// (6, 5, 'neigh_op_top_3')
// (6, 5, 'sp4_r_v_b_34')
// (6, 6, 'lutff_3/out')
// (6, 6, 'sp4_r_v_b_23')
// (6, 7, 'neigh_op_bot_3')
// (6, 7, 'sp4_r_v_b_10')
// (7, 0, 'span4_horz_l_12')
// (7, 0, 'span4_vert_25')
// (7, 1, 'sp4_v_b_25')
// (7, 2, 'sp4_v_b_12')
// (7, 3, 'sp4_v_b_1')
// (7, 3, 'sp4_v_t_47')
// (7, 4, 'sp4_v_b_47')
// (7, 5, 'neigh_op_tnl_3')
// (7, 5, 'sp4_v_b_34')
// (7, 6, 'neigh_op_lft_3')
// (7, 6, 'sp4_v_b_23')
// (7, 7, 'neigh_op_bnl_3')
// (7, 7, 'sp4_v_b_10')

wire n113;
// (3, 1, 'neigh_op_tnr_0')
// (3, 2, 'neigh_op_rgt_0')
// (3, 3, 'neigh_op_bnr_0')
// (4, 1, 'neigh_op_top_0')
// (4, 2, 'local_g3_0')
// (4, 2, 'lutff_0/out')
// (4, 2, 'lutff_1/in_2')
// (4, 2, 'lutff_7/in_0')
// (4, 3, 'neigh_op_bot_0')
// (5, 1, 'neigh_op_tnl_0')
// (5, 2, 'local_g0_0')
// (5, 2, 'lutff_6/in_0')
// (5, 2, 'neigh_op_lft_0')
// (5, 3, 'neigh_op_bnl_0')

wire n114;
// (3, 1, 'neigh_op_tnr_1')
// (3, 2, 'neigh_op_rgt_1')
// (3, 3, 'neigh_op_bnr_1')
// (4, 1, 'neigh_op_top_1')
// (4, 2, 'local_g2_1')
// (4, 2, 'lutff_1/out')
// (4, 2, 'lutff_4/in_3')
// (4, 3, 'neigh_op_bot_1')
// (5, 1, 'neigh_op_tnl_1')
// (5, 2, 'neigh_op_lft_1')
// (5, 3, 'neigh_op_bnl_1')

wire n115;
// (3, 1, 'neigh_op_tnr_2')
// (3, 2, 'neigh_op_rgt_2')
// (3, 3, 'neigh_op_bnr_2')
// (4, 0, 'span12_vert_23')
// (4, 1, 'neigh_op_top_2')
// (4, 1, 'sp12_v_b_23')
// (4, 2, 'lutff_2/out')
// (4, 2, 'sp12_v_b_20')
// (4, 3, 'local_g3_3')
// (4, 3, 'lutff_global/cen')
// (4, 3, 'neigh_op_bot_2')
// (4, 3, 'sp12_v_b_19')
// (4, 4, 'sp12_v_b_16')
// (4, 5, 'sp12_v_b_15')
// (4, 6, 'sp12_v_b_12')
// (4, 7, 'sp12_v_b_11')
// (4, 8, 'sp12_v_b_8')
// (4, 9, 'sp12_v_b_7')
// (4, 10, 'sp12_v_b_4')
// (4, 11, 'sp12_v_b_3')
// (4, 12, 'sp12_v_b_0')
// (5, 1, 'neigh_op_tnl_2')
// (5, 2, 'neigh_op_lft_2')
// (5, 3, 'neigh_op_bnl_2')

wire n116;
// (3, 1, 'neigh_op_tnr_3')
// (3, 2, 'neigh_op_rgt_3')
// (3, 3, 'neigh_op_bnr_3')
// (4, 1, 'neigh_op_top_3')
// (4, 2, 'lutff_3/out')
// (4, 3, 'neigh_op_bot_3')
// (5, 1, 'neigh_op_tnl_3')
// (5, 2, 'local_g1_3')
// (5, 2, 'lutff_2/in_2')
// (5, 2, 'lutff_4/in_2')
// (5, 2, 'neigh_op_lft_3')
// (5, 3, 'neigh_op_bnl_3')

wire n117;
// (3, 1, 'neigh_op_tnr_4')
// (3, 2, 'neigh_op_rgt_4')
// (3, 2, 'sp4_r_v_b_40')
// (3, 3, 'neigh_op_bnr_4')
// (3, 3, 'sp4_r_v_b_29')
// (3, 4, 'sp4_r_v_b_16')
// (3, 5, 'sp4_r_v_b_5')
// (4, 1, 'neigh_op_top_4')
// (4, 1, 'sp4_v_t_40')
// (4, 2, 'lutff_4/out')
// (4, 2, 'sp4_v_b_40')
// (4, 3, 'local_g0_4')
// (4, 3, 'local_g2_5')
// (4, 3, 'lutff_2/in_0')
// (4, 3, 'lutff_3/in_0')
// (4, 3, 'lutff_6/in_0')
// (4, 3, 'neigh_op_bot_4')
// (4, 3, 'sp4_v_b_29')
// (4, 4, 'sp4_v_b_16')
// (4, 5, 'sp4_v_b_5')
// (5, 1, 'neigh_op_tnl_4')
// (5, 2, 'neigh_op_lft_4')
// (5, 3, 'neigh_op_bnl_4')

wire n118;
// (3, 1, 'neigh_op_tnr_6')
// (3, 2, 'neigh_op_rgt_6')
// (3, 3, 'neigh_op_bnr_6')
// (4, 1, 'neigh_op_top_6')
// (4, 2, 'local_g3_6')
// (4, 2, 'lutff_4/in_1')
// (4, 2, 'lutff_6/out')
// (4, 3, 'neigh_op_bot_6')
// (5, 1, 'neigh_op_tnl_6')
// (5, 2, 'local_g0_6')
// (5, 2, 'lutff_3/in_1')
// (5, 2, 'lutff_4/in_0')
// (5, 2, 'lutff_5/in_1')
// (5, 2, 'neigh_op_lft_6')
// (5, 3, 'neigh_op_bnl_6')

wire \d_out[6] ;
// (3, 1, 'sp4_r_v_b_9')
// (3, 2, 'sp4_r_v_b_44')
// (3, 3, 'sp4_r_v_b_33')
// (3, 4, 'sp4_r_v_b_20')
// (3, 5, 'sp4_r_v_b_9')
// (4, 0, 'io_1/D_OUT_0')
// (4, 0, 'io_1/PAD')
// (4, 0, 'local_g0_1')
// (4, 0, 'span4_vert_9')
// (4, 1, 'sp4_v_b_9')
// (4, 1, 'sp4_v_t_44')
// (4, 2, 'sp4_v_b_44')
// (4, 3, 'sp4_v_b_33')
// (4, 4, 'neigh_op_tnr_2')
// (4, 4, 'sp4_v_b_20')
// (4, 5, 'neigh_op_rgt_2')
// (4, 5, 'sp4_h_r_9')
// (4, 5, 'sp4_v_b_9')
// (4, 6, 'neigh_op_bnr_2')
// (5, 4, 'neigh_op_top_2')
// (5, 5, 'lutff_2/out')
// (5, 5, 'sp4_h_r_20')
// (5, 6, 'neigh_op_bot_2')
// (6, 4, 'neigh_op_tnl_2')
// (6, 5, 'neigh_op_lft_2')
// (6, 5, 'sp4_h_r_33')
// (6, 6, 'neigh_op_bnl_2')
// (7, 5, 'sp4_h_r_44')
// (8, 5, 'sp4_h_l_44')

reg n120 = 0;
// (3, 2, 'neigh_op_tnr_2')
// (3, 3, 'neigh_op_rgt_2')
// (3, 4, 'neigh_op_bnr_2')
// (4, 2, 'local_g0_2')
// (4, 2, 'local_g1_2')
// (4, 2, 'lutff_0/in_1')
// (4, 2, 'lutff_3/in_1')
// (4, 2, 'lutff_5/in_1')
// (4, 2, 'lutff_6/in_1')
// (4, 2, 'neigh_op_top_2')
// (4, 3, 'local_g0_2')
// (4, 3, 'lutff_2/in_2')
// (4, 3, 'lutff_2/out')
// (4, 4, 'neigh_op_bot_2')
// (5, 2, 'neigh_op_tnl_2')
// (5, 3, 'neigh_op_lft_2')
// (5, 4, 'neigh_op_bnl_2')

reg n121 = 0;
// (3, 2, 'neigh_op_tnr_3')
// (3, 3, 'neigh_op_rgt_3')
// (3, 4, 'neigh_op_bnr_3')
// (4, 2, 'local_g0_3')
// (4, 2, 'local_g1_3')
// (4, 2, 'lutff_0/in_0')
// (4, 2, 'lutff_3/in_0')
// (4, 2, 'lutff_5/in_0')
// (4, 2, 'lutff_6/in_0')
// (4, 2, 'neigh_op_top_3')
// (4, 3, 'local_g0_3')
// (4, 3, 'lutff_3/in_2')
// (4, 3, 'lutff_3/out')
// (4, 4, 'neigh_op_bot_3')
// (5, 2, 'neigh_op_tnl_3')
// (5, 3, 'neigh_op_lft_3')
// (5, 4, 'neigh_op_bnl_3')

reg n122 = 0;
// (3, 2, 'neigh_op_tnr_4')
// (3, 3, 'neigh_op_rgt_4')
// (3, 4, 'neigh_op_bnr_4')
// (4, 2, 'local_g0_4')
// (4, 2, 'local_g1_4')
// (4, 2, 'lutff_0/in_3')
// (4, 2, 'lutff_3/in_3')
// (4, 2, 'lutff_5/in_3')
// (4, 2, 'lutff_6/in_3')
// (4, 2, 'neigh_op_top_4')
// (4, 3, 'local_g1_4')
// (4, 3, 'lutff_0/in_1')
// (4, 3, 'lutff_4/in_3')
// (4, 3, 'lutff_4/out')
// (4, 3, 'lutff_6/in_3')
// (4, 4, 'neigh_op_bot_4')
// (5, 2, 'neigh_op_tnl_4')
// (5, 3, 'neigh_op_lft_4')
// (5, 4, 'neigh_op_bnl_4')

reg n123 = 0;
// (3, 2, 'neigh_op_tnr_6')
// (3, 3, 'neigh_op_rgt_6')
// (3, 4, 'neigh_op_bnr_6')
// (4, 2, 'local_g0_6')
// (4, 2, 'local_g1_6')
// (4, 2, 'lutff_0/in_2')
// (4, 2, 'lutff_3/in_2')
// (4, 2, 'lutff_5/in_2')
// (4, 2, 'lutff_6/in_2')
// (4, 2, 'neigh_op_top_6')
// (4, 3, 'local_g0_6')
// (4, 3, 'local_g1_6')
// (4, 3, 'lutff_1/in_2')
// (4, 3, 'lutff_6/in_2')
// (4, 3, 'lutff_6/out')
// (4, 4, 'neigh_op_bot_6')
// (5, 2, 'neigh_op_tnl_6')
// (5, 3, 'neigh_op_lft_6')
// (5, 4, 'neigh_op_bnl_6')

wire \d_out[7] ;
// (3, 4, 'neigh_op_tnr_4')
// (3, 5, 'neigh_op_rgt_4')
// (3, 6, 'neigh_op_bnr_4')
// (4, 0, 'io_0/D_OUT_0')
// (4, 0, 'io_0/PAD')
// (4, 0, 'local_g0_0')
// (4, 0, 'span12_vert_16')
// (4, 1, 'sp12_v_b_16')
// (4, 2, 'sp12_v_b_15')
// (4, 3, 'sp12_v_b_12')
// (4, 4, 'neigh_op_top_4')
// (4, 4, 'sp12_v_b_11')
// (4, 5, 'lutff_4/out')
// (4, 5, 'sp12_v_b_8')
// (4, 6, 'neigh_op_bot_4')
// (4, 6, 'sp12_v_b_7')
// (4, 7, 'sp12_v_b_4')
// (4, 8, 'sp12_v_b_3')
// (4, 9, 'sp12_v_b_0')
// (5, 4, 'neigh_op_tnl_4')
// (5, 5, 'neigh_op_lft_4')
// (5, 6, 'neigh_op_bnl_4')

reg n125 = 0;
// (3, 4, 'neigh_op_tnr_5')
// (3, 5, 'neigh_op_rgt_5')
// (3, 6, 'neigh_op_bnr_5')
// (4, 4, 'neigh_op_top_5')
// (4, 5, 'local_g0_5')
// (4, 5, 'lutff_4/in_1')
// (4, 5, 'lutff_5/out')
// (4, 6, 'neigh_op_bot_5')
// (5, 4, 'neigh_op_tnl_5')
// (5, 5, 'neigh_op_lft_5')
// (5, 6, 'neigh_op_bnl_5')

wire n126;
// (3, 4, 'sp4_h_r_10')
// (4, 3, 'neigh_op_tnr_1')
// (4, 4, 'neigh_op_rgt_1')
// (4, 4, 'sp4_h_r_23')
// (4, 5, 'neigh_op_bnr_1')
// (5, 3, 'neigh_op_top_1')
// (5, 4, 'lutff_1/out')
// (5, 4, 'sp4_h_r_34')
// (5, 5, 'neigh_op_bot_1')
// (6, 3, 'neigh_op_tnl_1')
// (6, 4, 'neigh_op_lft_1')
// (6, 4, 'sp4_h_r_47')
// (6, 5, 'neigh_op_bnl_1')
// (7, 4, 'sp4_h_l_47')
// (7, 4, 'sp4_h_r_6')
// (8, 4, 'local_g0_3')
// (8, 4, 'lutff_2/in_3')
// (8, 4, 'lutff_6/in_3')
// (8, 4, 'sp4_h_r_19')
// (9, 4, 'sp4_h_r_30')
// (10, 4, 'sp4_h_r_43')
// (11, 4, 'sp4_h_l_43')

wire n127;
// (3, 4, 'sp4_r_v_b_39')
// (3, 5, 'sp4_r_v_b_26')
// (3, 6, 'sp4_r_v_b_15')
// (3, 7, 'sp4_r_v_b_2')
// (4, 3, 'sp4_v_t_39')
// (4, 4, 'sp4_v_b_39')
// (4, 5, 'sp4_v_b_26')
// (4, 6, 'local_g0_7')
// (4, 6, 'local_g2_2')
// (4, 6, 'lutff_1/in_3')
// (4, 6, 'lutff_6/in_3')
// (4, 6, 'neigh_op_tnr_2')
// (4, 6, 'sp4_v_b_15')
// (4, 7, 'local_g3_2')
// (4, 7, 'lutff_0/in_1')
// (4, 7, 'lutff_5/in_2')
// (4, 7, 'neigh_op_rgt_2')
// (4, 7, 'sp4_h_r_9')
// (4, 7, 'sp4_v_b_2')
// (4, 8, 'neigh_op_bnr_2')
// (5, 6, 'local_g1_2')
// (5, 6, 'lutff_6/in_1')
// (5, 6, 'neigh_op_top_2')
// (5, 7, 'lutff_2/out')
// (5, 7, 'sp4_h_r_20')
// (5, 8, 'neigh_op_bot_2')
// (6, 6, 'neigh_op_tnl_2')
// (6, 7, 'neigh_op_lft_2')
// (6, 7, 'sp4_h_r_33')
// (6, 8, 'neigh_op_bnl_2')
// (7, 7, 'sp4_h_r_44')
// (8, 7, 'sp4_h_l_44')

wire n128;
// (3, 5, 'neigh_op_tnr_0')
// (3, 6, 'neigh_op_rgt_0')
// (3, 7, 'neigh_op_bnr_0')
// (4, 4, 'sp4_r_v_b_41')
// (4, 5, 'neigh_op_top_0')
// (4, 5, 'sp4_r_v_b_28')
// (4, 6, 'lutff_0/out')
// (4, 6, 'sp4_r_v_b_17')
// (4, 7, 'local_g0_0')
// (4, 7, 'local_g1_0')
// (4, 7, 'lutff_6/in_3')
// (4, 7, 'lutff_7/in_1')
// (4, 7, 'neigh_op_bot_0')
// (4, 7, 'sp4_r_v_b_4')
// (5, 3, 'sp4_v_t_41')
// (5, 4, 'sp4_v_b_41')
// (5, 5, 'neigh_op_tnl_0')
// (5, 5, 'sp4_v_b_28')
// (5, 6, 'neigh_op_lft_0')
// (5, 6, 'sp4_v_b_17')
// (5, 7, 'local_g1_4')
// (5, 7, 'local_g2_0')
// (5, 7, 'lutff_3/in_1')
// (5, 7, 'lutff_7/in_0')
// (5, 7, 'neigh_op_bnl_0')
// (5, 7, 'sp4_h_r_4')
// (5, 7, 'sp4_v_b_4')
// (6, 7, 'local_g0_1')
// (6, 7, 'local_g1_1')
// (6, 7, 'lutff_0/in_2')
// (6, 7, 'lutff_1/in_0')
// (6, 7, 'lutff_4/in_2')
// (6, 7, 'lutff_6/in_2')
// (6, 7, 'sp4_h_r_17')
// (7, 7, 'sp4_h_r_28')
// (8, 7, 'sp4_h_r_41')
// (9, 7, 'sp4_h_l_41')

wire n129;
// (3, 5, 'neigh_op_tnr_1')
// (3, 6, 'neigh_op_rgt_1')
// (3, 7, 'neigh_op_bnr_1')
// (4, 5, 'neigh_op_top_1')
// (4, 6, 'local_g0_1')
// (4, 6, 'local_g1_1')
// (4, 6, 'lutff_0/in_2')
// (4, 6, 'lutff_1/out')
// (4, 6, 'lutff_2/in_1')
// (4, 6, 'lutff_3/in_2')
// (4, 7, 'neigh_op_bot_1')
// (5, 5, 'neigh_op_tnl_1')
// (5, 6, 'neigh_op_lft_1')
// (5, 7, 'neigh_op_bnl_1')

wire n130;
// (3, 5, 'neigh_op_tnr_2')
// (3, 6, 'neigh_op_rgt_2')
// (3, 7, 'neigh_op_bnr_2')
// (4, 4, 'sp4_r_v_b_45')
// (4, 5, 'neigh_op_top_2')
// (4, 5, 'sp4_r_v_b_32')
// (4, 6, 'lutff_2/out')
// (4, 6, 'sp4_r_v_b_21')
// (4, 7, 'local_g1_2')
// (4, 7, 'lutff_6/in_1')
// (4, 7, 'lutff_7/in_2')
// (4, 7, 'neigh_op_bot_2')
// (4, 7, 'sp4_r_v_b_8')
// (5, 3, 'sp4_v_t_45')
// (5, 4, 'sp4_v_b_45')
// (5, 5, 'neigh_op_tnl_2')
// (5, 5, 'sp4_v_b_32')
// (5, 6, 'neigh_op_lft_2')
// (5, 6, 'sp4_v_b_21')
// (5, 7, 'local_g2_2')
// (5, 7, 'local_g3_2')
// (5, 7, 'lutff_3/in_2')
// (5, 7, 'lutff_7/in_3')
// (5, 7, 'neigh_op_bnl_2')
// (5, 7, 'sp4_h_r_8')
// (5, 7, 'sp4_v_b_8')
// (6, 7, 'local_g0_5')
// (6, 7, 'local_g1_5')
// (6, 7, 'lutff_0/in_3')
// (6, 7, 'lutff_1/in_1')
// (6, 7, 'lutff_4/in_0')
// (6, 7, 'lutff_6/in_1')
// (6, 7, 'sp4_h_r_21')
// (7, 7, 'sp4_h_r_32')
// (8, 7, 'sp4_h_r_45')
// (9, 7, 'sp4_h_l_45')

wire n131;
// (3, 5, 'neigh_op_tnr_3')
// (3, 6, 'neigh_op_rgt_3')
// (3, 6, 'sp4_h_r_11')
// (3, 7, 'neigh_op_bnr_3')
// (4, 5, 'neigh_op_top_3')
// (4, 6, 'lutff_3/out')
// (4, 6, 'sp4_h_r_22')
// (4, 7, 'local_g0_3')
// (4, 7, 'local_g1_3')
// (4, 7, 'lutff_6/in_0')
// (4, 7, 'lutff_7/in_0')
// (4, 7, 'neigh_op_bot_3')
// (5, 5, 'neigh_op_tnl_3')
// (5, 6, 'neigh_op_lft_3')
// (5, 6, 'sp4_h_r_35')
// (5, 7, 'local_g2_3')
// (5, 7, 'lutff_3/in_0')
// (5, 7, 'lutff_7/in_2')
// (5, 7, 'neigh_op_bnl_3')
// (6, 6, 'sp4_h_r_46')
// (6, 7, 'local_g3_1')
// (6, 7, 'local_g3_6')
// (6, 7, 'lutff_0/in_0')
// (6, 7, 'lutff_1/in_2')
// (6, 7, 'lutff_4/in_3')
// (6, 7, 'lutff_6/in_3')
// (6, 7, 'sp4_r_v_b_41')
// (6, 7, 'sp4_r_v_b_46')
// (6, 8, 'sp4_r_v_b_28')
// (6, 8, 'sp4_r_v_b_35')
// (6, 9, 'sp4_r_v_b_17')
// (6, 9, 'sp4_r_v_b_22')
// (6, 10, 'sp4_r_v_b_11')
// (6, 10, 'sp4_r_v_b_4')
// (7, 6, 'sp4_h_l_46')
// (7, 6, 'sp4_v_t_41')
// (7, 6, 'sp4_v_t_46')
// (7, 7, 'sp4_v_b_41')
// (7, 7, 'sp4_v_b_46')
// (7, 8, 'sp4_v_b_28')
// (7, 8, 'sp4_v_b_35')
// (7, 9, 'sp4_v_b_17')
// (7, 9, 'sp4_v_b_22')
// (7, 10, 'sp4_v_b_11')
// (7, 10, 'sp4_v_b_4')

wire n132;
// (3, 6, 'neigh_op_tnr_0')
// (3, 7, 'neigh_op_rgt_0')
// (3, 8, 'neigh_op_bnr_0')
// (4, 3, 'sp12_v_t_23')
// (4, 4, 'sp12_v_b_23')
// (4, 5, 'sp12_v_b_20')
// (4, 6, 'neigh_op_top_0')
// (4, 6, 'sp12_v_b_19')
// (4, 7, 'lutff_0/out')
// (4, 7, 'sp12_v_b_16')
// (4, 8, 'local_g1_0')
// (4, 8, 'local_g3_7')
// (4, 8, 'lutff_0/in_2')
// (4, 8, 'lutff_4/in_1')
// (4, 8, 'lutff_5/in_1')
// (4, 8, 'lutff_6/in_2')
// (4, 8, 'neigh_op_bot_0')
// (4, 8, 'sp12_v_b_15')
// (4, 9, 'sp12_v_b_12')
// (4, 10, 'sp12_v_b_11')
// (4, 11, 'sp12_v_b_8')
// (4, 12, 'sp12_v_b_7')
// (4, 13, 'sp12_v_b_4')
// (4, 14, 'sp12_v_b_3')
// (4, 15, 'sp12_v_b_0')
// (5, 6, 'neigh_op_tnl_0')
// (5, 7, 'neigh_op_lft_0')
// (5, 8, 'neigh_op_bnl_0')

wire n133;
// (3, 6, 'neigh_op_tnr_2')
// (3, 7, 'neigh_op_rgt_2')
// (3, 8, 'neigh_op_bnr_2')
// (4, 5, 'sp4_r_v_b_45')
// (4, 6, 'neigh_op_top_2')
// (4, 6, 'sp4_r_v_b_32')
// (4, 7, 'lutff_2/out')
// (4, 7, 'sp4_r_v_b_21')
// (4, 7, 'sp4_r_v_b_37')
// (4, 8, 'local_g0_2')
// (4, 8, 'local_g1_2')
// (4, 8, 'lutff_4/in_0')
// (4, 8, 'lutff_5/in_0')
// (4, 8, 'lutff_7/in_2')
// (4, 8, 'neigh_op_bot_2')
// (4, 8, 'sp4_r_v_b_24')
// (4, 8, 'sp4_r_v_b_8')
// (4, 9, 'sp4_r_v_b_13')
// (4, 10, 'sp4_r_v_b_0')
// (5, 4, 'sp4_v_t_45')
// (5, 5, 'sp4_v_b_45')
// (5, 6, 'neigh_op_tnl_2')
// (5, 6, 'sp4_v_b_32')
// (5, 6, 'sp4_v_t_37')
// (5, 7, 'neigh_op_lft_2')
// (5, 7, 'sp4_v_b_21')
// (5, 7, 'sp4_v_b_37')
// (5, 8, 'local_g0_0')
// (5, 8, 'lutff_4/in_0')
// (5, 8, 'neigh_op_bnl_2')
// (5, 8, 'sp4_v_b_24')
// (5, 8, 'sp4_v_b_8')
// (5, 9, 'local_g0_5')
// (5, 9, 'lutff_5/in_2')
// (5, 9, 'sp4_v_b_13')
// (5, 10, 'sp4_v_b_0')

wire n134;
// (3, 6, 'neigh_op_tnr_5')
// (3, 7, 'neigh_op_rgt_5')
// (3, 8, 'neigh_op_bnr_5')
// (4, 6, 'neigh_op_top_5')
// (4, 7, 'lutff_5/out')
// (4, 8, 'local_g1_5')
// (4, 8, 'lutff_3/in_3')
// (4, 8, 'neigh_op_bot_5')
// (5, 6, 'neigh_op_tnl_5')
// (5, 7, 'neigh_op_lft_5')
// (5, 8, 'local_g3_5')
// (5, 8, 'lutff_5/in_1')
// (5, 8, 'neigh_op_bnl_5')

wire n135;
// (3, 6, 'neigh_op_tnr_6')
// (3, 7, 'neigh_op_rgt_6')
// (3, 8, 'neigh_op_bnr_6')
// (4, 6, 'neigh_op_top_6')
// (4, 7, 'local_g0_6')
// (4, 7, 'local_g1_6')
// (4, 7, 'lutff_0/in_2')
// (4, 7, 'lutff_1/in_1')
// (4, 7, 'lutff_2/in_1')
// (4, 7, 'lutff_5/in_1')
// (4, 7, 'lutff_6/out')
// (4, 8, 'neigh_op_bot_6')
// (5, 6, 'neigh_op_tnl_6')
// (5, 7, 'neigh_op_lft_6')
// (5, 8, 'neigh_op_bnl_6')

wire n136;
// (3, 6, 'neigh_op_tnr_7')
// (3, 7, 'neigh_op_rgt_7')
// (3, 8, 'neigh_op_bnr_7')
// (4, 6, 'neigh_op_top_7')
// (4, 7, 'local_g2_7')
// (4, 7, 'local_g3_7')
// (4, 7, 'lutff_0/in_0')
// (4, 7, 'lutff_1/in_0')
// (4, 7, 'lutff_2/in_0')
// (4, 7, 'lutff_5/in_0')
// (4, 7, 'lutff_7/out')
// (4, 8, 'neigh_op_bot_7')
// (5, 6, 'neigh_op_tnl_7')
// (5, 7, 'neigh_op_lft_7')
// (5, 8, 'neigh_op_bnl_7')

reg n137 = 0;
// (3, 6, 'sp12_h_r_0')
// (4, 6, 'sp12_h_r_3')
// (5, 6, 'sp12_h_r_4')
// (5, 7, 'sp4_r_v_b_40')
// (5, 8, 'sp4_r_v_b_29')
// (5, 9, 'sp4_r_v_b_16')
// (5, 10, 'sp4_r_v_b_5')
// (5, 11, 'sp4_r_v_b_40')
// (5, 11, 'sp4_r_v_b_45')
// (5, 12, 'sp4_r_v_b_29')
// (5, 12, 'sp4_r_v_b_32')
// (5, 13, 'sp4_r_v_b_16')
// (5, 13, 'sp4_r_v_b_21')
// (5, 14, 'sp4_r_v_b_5')
// (5, 14, 'sp4_r_v_b_8')
// (6, 6, 'sp12_h_r_7')
// (6, 6, 'sp4_h_r_5')
// (6, 6, 'sp4_v_t_40')
// (6, 7, 'sp4_v_b_40')
// (6, 8, 'sp4_v_b_29')
// (6, 9, 'sp4_v_b_16')
// (6, 10, 'sp4_v_b_5')
// (6, 10, 'sp4_v_t_40')
// (6, 10, 'sp4_v_t_45')
// (6, 11, 'sp4_v_b_40')
// (6, 11, 'sp4_v_b_45')
// (6, 12, 'sp4_v_b_29')
// (6, 12, 'sp4_v_b_32')
// (6, 13, 'local_g0_0')
// (6, 13, 'local_g0_5')
// (6, 13, 'lutff_0/in_2')
// (6, 13, 'lutff_3/in_2')
// (6, 13, 'sp4_v_b_16')
// (6, 13, 'sp4_v_b_21')
// (6, 14, 'sp4_v_b_5')
// (6, 14, 'sp4_v_b_8')
// (7, 6, 'sp12_h_r_8')
// (7, 6, 'sp4_h_r_16')
// (8, 5, 'neigh_op_tnr_2')
// (8, 6, 'neigh_op_rgt_2')
// (8, 6, 'sp12_h_r_11')
// (8, 6, 'sp4_h_r_29')
// (8, 7, 'neigh_op_bnr_2')
// (8, 11, 'sp4_r_v_b_39')
// (8, 12, 'local_g0_2')
// (8, 12, 'lutff_4/in_0')
// (8, 12, 'sp4_r_v_b_26')
// (8, 13, 'sp4_r_v_b_15')
// (8, 14, 'sp4_r_v_b_2')
// (9, 4, 'sp12_v_t_23')
// (9, 5, 'neigh_op_top_2')
// (9, 5, 'sp12_v_b_23')
// (9, 6, 'lutff_2/out')
// (9, 6, 'sp12_h_r_12')
// (9, 6, 'sp12_v_b_20')
// (9, 6, 'sp4_h_r_40')
// (9, 7, 'neigh_op_bot_2')
// (9, 7, 'sp12_v_b_19')
// (9, 8, 'sp12_v_b_16')
// (9, 9, 'sp12_v_b_15')
// (9, 10, 'sp12_v_b_12')
// (9, 10, 'sp4_v_t_39')
// (9, 11, 'sp12_v_b_11')
// (9, 11, 'sp4_v_b_39')
// (9, 12, 'sp12_v_b_8')
// (9, 12, 'sp4_v_b_26')
// (9, 13, 'sp12_v_b_7')
// (9, 13, 'sp4_v_b_15')
// (9, 14, 'sp12_v_b_4')
// (9, 14, 'sp4_v_b_2')
// (9, 15, 'sp12_v_b_3')
// (9, 16, 'sp12_v_b_0')
// (10, 5, 'neigh_op_tnl_2')
// (10, 6, 'neigh_op_lft_2')
// (10, 6, 'sp12_h_r_15')
// (10, 6, 'sp4_h_l_40')
// (10, 7, 'neigh_op_bnl_2')
// (11, 6, 'local_g0_0')
// (11, 6, 'lutff_2/in_0')
// (11, 6, 'sp12_h_r_16')
// (12, 6, 'sp12_h_r_19')
// (13, 6, 'span12_horz_19')

wire n138;
// (3, 7, 'neigh_op_tnr_0')
// (3, 7, 'sp4_r_v_b_45')
// (3, 8, 'neigh_op_rgt_0')
// (3, 8, 'sp4_r_v_b_32')
// (3, 9, 'neigh_op_bnr_0')
// (3, 9, 'sp4_r_v_b_21')
// (3, 10, 'sp4_r_v_b_8')
// (4, 6, 'sp4_v_t_45')
// (4, 7, 'neigh_op_top_0')
// (4, 7, 'sp4_v_b_45')
// (4, 8, 'local_g0_0')
// (4, 8, 'lutff_0/out')
// (4, 8, 'lutff_3/in_1')
// (4, 8, 'sp4_v_b_32')
// (4, 9, 'local_g1_0')
// (4, 9, 'lutff_1/in_2')
// (4, 9, 'neigh_op_bot_0')
// (4, 9, 'sp4_v_b_21')
// (4, 10, 'local_g1_0')
// (4, 10, 'lutff_2/in_3')
// (4, 10, 'sp4_v_b_8')
// (5, 7, 'neigh_op_tnl_0')
// (5, 8, 'neigh_op_lft_0')
// (5, 9, 'neigh_op_bnl_0')

wire n139;
// (3, 7, 'neigh_op_tnr_2')
// (3, 8, 'neigh_op_rgt_2')
// (3, 9, 'neigh_op_bnr_2')
// (4, 7, 'neigh_op_top_2')
// (4, 8, 'lutff_2/out')
// (4, 9, 'local_g0_2')
// (4, 9, 'lutff_5/in_3')
// (4, 9, 'neigh_op_bot_2')
// (5, 7, 'neigh_op_tnl_2')
// (5, 8, 'neigh_op_lft_2')
// (5, 9, 'neigh_op_bnl_2')

wire n140;
// (3, 7, 'neigh_op_tnr_3')
// (3, 8, 'neigh_op_rgt_3')
// (3, 9, 'neigh_op_bnr_3')
// (4, 7, 'neigh_op_top_3')
// (4, 8, 'lutff_3/out')
// (4, 8, 'sp4_h_r_6')
// (4, 8, 'sp4_r_v_b_39')
// (4, 9, 'neigh_op_bot_3')
// (4, 9, 'sp4_r_v_b_26')
// (4, 10, 'sp4_r_v_b_15')
// (4, 11, 'sp4_r_v_b_2')
// (5, 7, 'neigh_op_tnl_3')
// (5, 7, 'sp4_v_t_39')
// (5, 8, 'neigh_op_lft_3')
// (5, 8, 'sp4_h_r_19')
// (5, 8, 'sp4_v_b_39')
// (5, 9, 'neigh_op_bnl_3')
// (5, 9, 'sp4_v_b_26')
// (5, 10, 'sp4_v_b_15')
// (5, 11, 'sp4_h_r_8')
// (5, 11, 'sp4_v_b_2')
// (6, 8, 'sp4_h_r_30')
// (6, 11, 'local_g0_5')
// (6, 11, 'lutff_4/in_3')
// (6, 11, 'lutff_7/in_2')
// (6, 11, 'sp4_h_r_21')
// (7, 8, 'sp4_h_r_43')
// (7, 9, 'sp4_r_v_b_43')
// (7, 10, 'local_g0_6')
// (7, 10, 'local_g1_6')
// (7, 10, 'lutff_2/in_3')
// (7, 10, 'lutff_3/in_3')
// (7, 10, 'lutff_6/in_2')
// (7, 10, 'sp4_r_v_b_30')
// (7, 11, 'sp4_h_r_32')
// (7, 11, 'sp4_r_v_b_19')
// (7, 12, 'sp4_r_v_b_6')
// (8, 8, 'sp4_h_l_43')
// (8, 8, 'sp4_v_t_43')
// (8, 9, 'sp4_v_b_43')
// (8, 10, 'sp4_v_b_30')
// (8, 11, 'sp4_h_r_45')
// (8, 11, 'sp4_v_b_19')
// (8, 12, 'sp4_v_b_6')
// (9, 11, 'sp4_h_l_45')
// (9, 11, 'sp4_h_r_11')
// (10, 11, 'sp4_h_r_22')
// (11, 11, 'local_g2_3')
// (11, 11, 'lutff_4/in_3')
// (11, 11, 'sp4_h_r_35')
// (12, 11, 'sp4_h_r_46')
// (13, 11, 'span4_horz_46')

wire n141;
// (3, 7, 'neigh_op_tnr_7')
// (3, 8, 'neigh_op_rgt_7')
// (3, 9, 'neigh_op_bnr_7')
// (4, 7, 'neigh_op_top_7')
// (4, 8, 'local_g0_7')
// (4, 8, 'lutff_3/in_0')
// (4, 8, 'lutff_7/out')
// (4, 9, 'neigh_op_bot_7')
// (5, 7, 'neigh_op_tnl_7')
// (5, 8, 'neigh_op_lft_7')
// (5, 9, 'neigh_op_bnl_7')

wire n142;
// (3, 7, 'sp12_h_r_0')
// (4, 7, 'sp12_h_r_3')
// (5, 7, 'sp12_h_r_4')
// (6, 6, 'neigh_op_tnr_0')
// (6, 7, 'neigh_op_rgt_0')
// (6, 7, 'sp12_h_r_7')
// (6, 8, 'neigh_op_bnr_0')
// (7, 5, 'sp4_r_v_b_41')
// (7, 6, 'neigh_op_top_0')
// (7, 6, 'sp4_r_v_b_28')
// (7, 7, 'lutff_0/out')
// (7, 7, 'sp12_h_r_8')
// (7, 7, 'sp4_r_v_b_17')
// (7, 8, 'neigh_op_bot_0')
// (7, 8, 'sp4_r_v_b_4')
// (8, 4, 'sp4_v_t_41')
// (8, 5, 'sp4_v_b_41')
// (8, 6, 'neigh_op_tnl_0')
// (8, 6, 'sp4_v_b_28')
// (8, 7, 'neigh_op_lft_0')
// (8, 7, 'sp12_h_r_11')
// (8, 7, 'sp4_h_r_7')
// (8, 7, 'sp4_v_b_17')
// (8, 8, 'neigh_op_bnl_0')
// (8, 8, 'sp4_h_r_10')
// (8, 8, 'sp4_v_b_4')
// (9, 7, 'local_g0_4')
// (9, 7, 'lutff_0/in_2')
// (9, 7, 'sp12_h_r_12')
// (9, 7, 'sp4_h_r_18')
// (9, 8, 'local_g0_7')
// (9, 8, 'lutff_5/in_0')
// (9, 8, 'sp4_h_r_23')
// (10, 7, 'sp12_h_r_15')
// (10, 7, 'sp4_h_r_31')
// (10, 8, 'sp4_h_r_34')
// (11, 7, 'sp12_h_r_16')
// (11, 7, 'sp4_h_r_42')
// (11, 8, 'sp4_h_r_47')
// (11, 8, 'sp4_r_v_b_42')
// (11, 9, 'local_g0_7')
// (11, 9, 'local_g2_6')
// (11, 9, 'lutff_1/in_2')
// (11, 9, 'lutff_6/in_2')
// (11, 9, 'sp4_r_v_b_31')
// (11, 9, 'sp4_r_v_b_38')
// (11, 10, 'sp4_r_v_b_18')
// (11, 10, 'sp4_r_v_b_27')
// (11, 11, 'sp4_r_v_b_14')
// (11, 11, 'sp4_r_v_b_7')
// (11, 12, 'sp4_r_v_b_3')
// (12, 7, 'sp12_h_r_19')
// (12, 7, 'sp4_h_l_42')
// (12, 7, 'sp4_v_t_42')
// (12, 8, 'sp4_h_l_47')
// (12, 8, 'sp4_v_b_42')
// (12, 8, 'sp4_v_t_38')
// (12, 9, 'sp4_v_b_31')
// (12, 9, 'sp4_v_b_38')
// (12, 10, 'sp4_v_b_18')
// (12, 10, 'sp4_v_b_27')
// (12, 11, 'sp4_v_b_14')
// (12, 11, 'sp4_v_b_7')
// (12, 12, 'sp4_v_b_3')
// (13, 7, 'span12_horz_19')

reg n143 = 0;
// (3, 7, 'sp12_h_r_1')
// (4, 7, 'sp12_h_r_2')
// (5, 6, 'neigh_op_tnr_7')
// (5, 7, 'neigh_op_rgt_7')
// (5, 7, 'sp12_h_r_5')
// (5, 8, 'neigh_op_bnr_7')
// (6, 6, 'neigh_op_top_7')
// (6, 7, 'lutff_7/out')
// (6, 7, 'sp12_h_r_6')
// (6, 8, 'neigh_op_bot_7')
// (7, 6, 'neigh_op_tnl_7')
// (7, 7, 'local_g0_1')
// (7, 7, 'lutff_5/in_0')
// (7, 7, 'neigh_op_lft_7')
// (7, 7, 'sp12_h_r_9')
// (7, 8, 'neigh_op_bnl_7')
// (8, 7, 'sp12_h_r_10')
// (9, 7, 'sp12_h_r_13')
// (10, 7, 'sp12_h_r_14')
// (11, 7, 'sp12_h_r_17')
// (12, 7, 'sp12_h_r_18')
// (13, 7, 'span12_horz_18')

wire n144;
// (3, 7, 'sp4_h_r_1')
// (4, 7, 'sp4_h_r_12')
// (5, 6, 'local_g2_2')
// (5, 6, 'local_g3_2')
// (5, 6, 'lutff_5/in_0')
// (5, 6, 'lutff_6/in_0')
// (5, 6, 'neigh_op_tnr_2')
// (5, 7, 'local_g2_1')
// (5, 7, 'lutff_4/in_3')
// (5, 7, 'neigh_op_rgt_2')
// (5, 7, 'sp4_h_r_25')
// (5, 8, 'neigh_op_bnr_2')
// (6, 6, 'neigh_op_top_2')
// (6, 7, 'local_g0_2')
// (6, 7, 'lutff_2/out')
// (6, 7, 'lutff_3/in_1')
// (6, 7, 'sp4_h_r_36')
// (6, 8, 'neigh_op_bot_2')
// (7, 6, 'neigh_op_tnl_2')
// (7, 7, 'neigh_op_lft_2')
// (7, 7, 'sp4_h_l_36')
// (7, 8, 'neigh_op_bnl_2')

reg n145 = 0;
// (3, 8, 'neigh_op_tnr_3')
// (3, 9, 'neigh_op_rgt_3')
// (3, 10, 'neigh_op_bnr_3')
// (4, 8, 'neigh_op_top_3')
// (4, 9, 'local_g0_3')
// (4, 9, 'lutff_2/in_1')
// (4, 9, 'lutff_3/out')
// (4, 10, 'local_g0_3')
// (4, 10, 'lutff_1/in_2')
// (4, 10, 'neigh_op_bot_3')
// (5, 8, 'neigh_op_tnl_3')
// (5, 9, 'neigh_op_lft_3')
// (5, 10, 'neigh_op_bnl_3')

wire n146;
// (3, 9, 'neigh_op_tnr_0')
// (3, 10, 'neigh_op_rgt_0')
// (3, 11, 'neigh_op_bnr_0')
// (4, 9, 'neigh_op_top_0')
// (4, 10, 'local_g0_0')
// (4, 10, 'local_g2_0')
// (4, 10, 'lutff_0/out')
// (4, 10, 'lutff_2/in_2')
// (4, 10, 'lutff_5/in_3')
// (4, 11, 'neigh_op_bot_0')
// (5, 9, 'neigh_op_tnl_0')
// (5, 10, 'neigh_op_lft_0')
// (5, 11, 'neigh_op_bnl_0')

wire n147;
// (3, 9, 'neigh_op_tnr_1')
// (3, 10, 'neigh_op_rgt_1')
// (3, 11, 'neigh_op_bnr_1')
// (4, 9, 'neigh_op_top_1')
// (4, 9, 'sp4_r_v_b_46')
// (4, 10, 'lutff_1/out')
// (4, 10, 'sp4_r_v_b_35')
// (4, 11, 'neigh_op_bot_1')
// (4, 11, 'sp4_r_v_b_22')
// (4, 12, 'sp4_r_v_b_11')
// (5, 8, 'sp4_v_t_46')
// (5, 9, 'neigh_op_tnl_1')
// (5, 9, 'sp4_v_b_46')
// (5, 10, 'neigh_op_lft_1')
// (5, 10, 'sp4_v_b_35')
// (5, 11, 'local_g2_1')
// (5, 11, 'lutff_2/in_1')
// (5, 11, 'neigh_op_bnl_1')
// (5, 11, 'sp4_v_b_22')
// (5, 12, 'local_g0_3')
// (5, 12, 'lutff_6/in_1')
// (5, 12, 'sp4_v_b_11')

reg n148 = 0;
// (3, 9, 'neigh_op_tnr_3')
// (3, 10, 'neigh_op_rgt_3')
// (3, 11, 'neigh_op_bnr_3')
// (4, 9, 'local_g1_3')
// (4, 9, 'lutff_3/in_1')
// (4, 9, 'neigh_op_top_3')
// (4, 10, 'local_g1_3')
// (4, 10, 'lutff_3/out')
// (4, 10, 'lutff_6/in_2')
// (4, 11, 'neigh_op_bot_3')
// (5, 9, 'neigh_op_tnl_3')
// (5, 10, 'neigh_op_lft_3')
// (5, 11, 'neigh_op_bnl_3')

reg n149 = 0;
// (3, 9, 'neigh_op_tnr_4')
// (3, 10, 'neigh_op_rgt_4')
// (3, 11, 'neigh_op_bnr_4')
// (4, 9, 'neigh_op_top_4')
// (4, 10, 'local_g3_4')
// (4, 10, 'lutff_4/out')
// (4, 10, 'lutff_5/in_2')
// (4, 11, 'neigh_op_bot_4')
// (5, 9, 'neigh_op_tnl_4')
// (5, 10, 'local_g1_4')
// (5, 10, 'lutff_1/in_0')
// (5, 10, 'neigh_op_lft_4')
// (5, 11, 'neigh_op_bnl_4')

reg n150 = 0;
// (3, 9, 'neigh_op_tnr_5')
// (3, 10, 'neigh_op_rgt_5')
// (3, 11, 'neigh_op_bnr_5')
// (4, 9, 'neigh_op_top_5')
// (4, 10, 'lutff_5/out')
// (4, 11, 'local_g1_5')
// (4, 11, 'lutff_2/in_2')
// (4, 11, 'lutff_3/in_1')
// (4, 11, 'neigh_op_bot_5')
// (5, 9, 'neigh_op_tnl_5')
// (5, 10, 'neigh_op_lft_5')
// (5, 11, 'neigh_op_bnl_5')

reg n151 = 0;
// (3, 9, 'neigh_op_tnr_6')
// (3, 10, 'neigh_op_rgt_6')
// (3, 11, 'neigh_op_bnr_6')
// (4, 9, 'neigh_op_top_6')
// (4, 10, 'local_g0_6')
// (4, 10, 'lutff_1/in_1')
// (4, 10, 'lutff_6/out')
// (4, 11, 'neigh_op_bot_6')
// (5, 9, 'neigh_op_tnl_6')
// (5, 10, 'neigh_op_lft_6')
// (5, 11, 'neigh_op_bnl_6')

reg n152 = 0;
// (3, 9, 'neigh_op_tnr_7')
// (3, 10, 'neigh_op_rgt_7')
// (3, 11, 'neigh_op_bnr_7')
// (4, 9, 'neigh_op_top_7')
// (4, 10, 'local_g0_7')
// (4, 10, 'lutff_6/in_1')
// (4, 10, 'lutff_7/out')
// (4, 11, 'neigh_op_bot_7')
// (5, 9, 'neigh_op_tnl_7')
// (5, 10, 'neigh_op_lft_7')
// (5, 11, 'neigh_op_bnl_7')

wire n153;
// (3, 10, 'neigh_op_tnr_1')
// (3, 11, 'neigh_op_rgt_1')
// (3, 12, 'neigh_op_bnr_1')
// (4, 10, 'neigh_op_top_1')
// (4, 11, 'lutff_1/out')
// (4, 12, 'neigh_op_bot_1')
// (5, 10, 'neigh_op_tnl_1')
// (5, 11, 'neigh_op_lft_1')
// (5, 12, 'local_g2_1')
// (5, 12, 'local_g3_1')
// (5, 12, 'lutff_0/in_1')
// (5, 12, 'lutff_7/in_1')
// (5, 12, 'neigh_op_bnl_1')

reg n154 = 0;
// (3, 10, 'neigh_op_tnr_2')
// (3, 11, 'neigh_op_rgt_2')
// (3, 12, 'neigh_op_bnr_2')
// (4, 10, 'neigh_op_top_2')
// (4, 11, 'local_g1_2')
// (4, 11, 'lutff_2/out')
// (4, 11, 'lutff_4/in_1')
// (4, 12, 'neigh_op_bot_2')
// (5, 10, 'neigh_op_tnl_2')
// (5, 11, 'neigh_op_lft_2')
// (5, 12, 'neigh_op_bnl_2')

reg n155 = 0;
// (3, 10, 'neigh_op_tnr_3')
// (3, 11, 'neigh_op_rgt_3')
// (3, 12, 'neigh_op_bnr_3')
// (4, 10, 'neigh_op_top_3')
// (4, 11, 'local_g1_3')
// (4, 11, 'lutff_3/out')
// (4, 11, 'lutff_4/in_2')
// (4, 11, 'lutff_5/in_1')
// (4, 12, 'neigh_op_bot_3')
// (5, 10, 'neigh_op_tnl_3')
// (5, 11, 'neigh_op_lft_3')
// (5, 12, 'neigh_op_bnl_3')

reg n156 = 0;
// (3, 10, 'neigh_op_tnr_4')
// (3, 11, 'neigh_op_rgt_4')
// (3, 12, 'neigh_op_bnr_4')
// (4, 10, 'neigh_op_top_4')
// (4, 11, 'local_g0_4')
// (4, 11, 'lutff_1/in_1')
// (4, 11, 'lutff_4/out')
// (4, 12, 'neigh_op_bot_4')
// (5, 10, 'neigh_op_tnl_4')
// (5, 11, 'neigh_op_lft_4')
// (5, 12, 'neigh_op_bnl_4')

reg n157 = 0;
// (3, 10, 'neigh_op_tnr_5')
// (3, 11, 'neigh_op_rgt_5')
// (3, 12, 'neigh_op_bnr_5')
// (4, 10, 'local_g0_5')
// (4, 10, 'lutff_4/in_1')
// (4, 10, 'neigh_op_top_5')
// (4, 11, 'local_g0_5')
// (4, 11, 'lutff_1/in_2')
// (4, 11, 'lutff_5/out')
// (4, 12, 'neigh_op_bot_5')
// (5, 10, 'neigh_op_tnl_5')
// (5, 11, 'neigh_op_lft_5')
// (5, 12, 'neigh_op_bnl_5')

reg n158 = 0;
// (3, 11, 'neigh_op_tnr_1')
// (3, 12, 'neigh_op_rgt_1')
// (3, 13, 'neigh_op_bnr_1')
// (4, 11, 'neigh_op_top_1')
// (4, 12, 'lutff_1/out')
// (4, 13, 'neigh_op_bot_1')
// (5, 11, 'neigh_op_tnl_1')
// (5, 12, 'local_g0_1')
// (5, 12, 'lutff_5/in_0')
// (5, 12, 'neigh_op_lft_1')
// (5, 13, 'neigh_op_bnl_1')

reg n159 = 0;
// (3, 11, 'neigh_op_tnr_3')
// (3, 12, 'neigh_op_rgt_3')
// (3, 13, 'neigh_op_bnr_3')
// (4, 11, 'neigh_op_top_3')
// (4, 12, 'local_g1_3')
// (4, 12, 'lutff_3/out')
// (4, 12, 'lutff_6/in_0')
// (4, 13, 'neigh_op_bot_3')
// (5, 11, 'neigh_op_tnl_3')
// (5, 12, 'neigh_op_lft_3')
// (5, 13, 'neigh_op_bnl_3')

reg n160 = 0;
// (3, 11, 'neigh_op_tnr_6')
// (3, 12, 'neigh_op_rgt_6')
// (3, 13, 'neigh_op_bnr_6')
// (4, 11, 'neigh_op_top_6')
// (4, 12, 'local_g0_6')
// (4, 12, 'lutff_4/in_0')
// (4, 12, 'lutff_6/out')
// (4, 13, 'neigh_op_bot_6')
// (5, 11, 'neigh_op_tnl_6')
// (5, 12, 'neigh_op_lft_6')
// (5, 13, 'neigh_op_bnl_6')

reg n161 = 0;
// (3, 11, 'neigh_op_tnr_7')
// (3, 12, 'neigh_op_rgt_7')
// (3, 13, 'neigh_op_bnr_7')
// (4, 11, 'neigh_op_top_7')
// (4, 12, 'lutff_7/out')
// (4, 13, 'local_g1_7')
// (4, 13, 'lutff_4/in_0')
// (4, 13, 'neigh_op_bot_7')
// (5, 11, 'neigh_op_tnl_7')
// (5, 12, 'neigh_op_lft_7')
// (5, 13, 'neigh_op_bnl_7')

wire n162;
// (3, 12, 'neigh_op_tnr_0')
// (3, 13, 'neigh_op_rgt_0')
// (3, 14, 'neigh_op_bnr_0')
// (4, 12, 'neigh_op_top_0')
// (4, 13, 'lutff_0/out')
// (4, 14, 'neigh_op_bot_0')
// (5, 12, 'local_g2_0')
// (5, 12, 'lutff_1/in_3')
// (5, 12, 'neigh_op_tnl_0')
// (5, 13, 'neigh_op_lft_0')
// (5, 14, 'neigh_op_bnl_0')

reg n163 = 0;
// (3, 12, 'neigh_op_tnr_3')
// (3, 13, 'neigh_op_rgt_3')
// (3, 14, 'neigh_op_bnr_3')
// (4, 12, 'neigh_op_top_3')
// (4, 13, 'local_g0_3')
// (4, 13, 'lutff_3/out')
// (4, 13, 'lutff_7/in_0')
// (4, 14, 'neigh_op_bot_3')
// (5, 12, 'neigh_op_tnl_3')
// (5, 13, 'neigh_op_lft_3')
// (5, 14, 'neigh_op_bnl_3')

reg n164 = 0;
// (3, 12, 'neigh_op_tnr_5')
// (3, 13, 'neigh_op_rgt_5')
// (3, 14, 'neigh_op_bnr_5')
// (4, 12, 'neigh_op_top_5')
// (4, 13, 'local_g1_5')
// (4, 13, 'lutff_5/out')
// (4, 13, 'lutff_6/in_0')
// (4, 14, 'neigh_op_bot_5')
// (5, 12, 'neigh_op_tnl_5')
// (5, 13, 'neigh_op_lft_5')
// (5, 14, 'neigh_op_bnl_5')

reg n165 = 0;
// (3, 12, 'neigh_op_tnr_6')
// (3, 13, 'neigh_op_rgt_6')
// (3, 14, 'neigh_op_bnr_6')
// (4, 12, 'neigh_op_top_6')
// (4, 13, 'local_g1_6')
// (4, 13, 'lutff_3/in_0')
// (4, 13, 'lutff_6/out')
// (4, 14, 'neigh_op_bot_6')
// (5, 12, 'neigh_op_tnl_6')
// (5, 13, 'neigh_op_lft_6')
// (5, 14, 'neigh_op_bnl_6')

wire n166;
// (4, 1, 'neigh_op_tnr_2')
// (4, 2, 'local_g2_2')
// (4, 2, 'lutff_4/in_2')
// (4, 2, 'neigh_op_rgt_2')
// (4, 3, 'neigh_op_bnr_2')
// (5, 1, 'neigh_op_top_2')
// (5, 2, 'local_g0_2')
// (5, 2, 'lutff_2/out')
// (5, 2, 'lutff_6/in_2')
// (5, 3, 'neigh_op_bot_2')
// (6, 1, 'neigh_op_tnl_2')
// (6, 2, 'neigh_op_lft_2')
// (6, 3, 'neigh_op_bnl_2')

wire n167;
// (4, 1, 'neigh_op_tnr_4')
// (4, 2, 'neigh_op_rgt_4')
// (4, 3, 'neigh_op_bnr_4')
// (5, 1, 'neigh_op_top_4')
// (5, 2, 'local_g1_4')
// (5, 2, 'lutff_4/out')
// (5, 2, 'lutff_7/in_2')
// (5, 3, 'neigh_op_bot_4')
// (6, 1, 'neigh_op_tnl_4')
// (6, 2, 'neigh_op_lft_4')
// (6, 3, 'neigh_op_bnl_4')

wire n168;
// (4, 1, 'sp4_r_v_b_41')
// (4, 2, 'sp4_r_v_b_28')
// (4, 3, 'local_g3_1')
// (4, 3, 'lutff_4/in_2')
// (4, 3, 'sp4_r_v_b_17')
// (4, 4, 'sp4_r_v_b_4')
// (5, 0, 'span4_vert_41')
// (5, 1, 'sp4_v_b_41')
// (5, 2, 'sp4_v_b_28')
// (5, 3, 'neigh_op_tnr_3')
// (5, 3, 'sp4_v_b_17')
// (5, 4, 'neigh_op_rgt_3')
// (5, 4, 'sp4_h_r_11')
// (5, 4, 'sp4_v_b_4')
// (5, 5, 'neigh_op_bnr_3')
// (6, 3, 'neigh_op_top_3')
// (6, 4, 'lutff_3/out')
// (6, 4, 'sp4_h_r_22')
// (6, 5, 'local_g0_3')
// (6, 5, 'lutff_1/in_0')
// (6, 5, 'neigh_op_bot_3')
// (7, 3, 'neigh_op_tnl_3')
// (7, 4, 'local_g0_3')
// (7, 4, 'lutff_4/in_3')
// (7, 4, 'lutff_6/in_3')
// (7, 4, 'neigh_op_lft_3')
// (7, 4, 'sp4_h_r_35')
// (7, 5, 'local_g2_3')
// (7, 5, 'local_g3_3')
// (7, 5, 'lutff_2/in_0')
// (7, 5, 'lutff_5/in_0')
// (7, 5, 'neigh_op_bnl_3')
// (8, 4, 'local_g3_6')
// (8, 4, 'lutff_7/in_0')
// (8, 4, 'sp4_h_r_46')
// (8, 5, 'local_g3_1')
// (8, 5, 'lutff_0/in_0')
// (8, 5, 'lutff_2/in_0')
// (8, 5, 'sp4_r_v_b_41')
// (8, 6, 'sp4_r_v_b_28')
// (8, 7, 'sp4_r_v_b_17')
// (8, 8, 'sp4_r_v_b_4')
// (9, 4, 'sp4_h_l_46')
// (9, 4, 'sp4_v_t_41')
// (9, 5, 'sp4_v_b_41')
// (9, 6, 'sp4_v_b_28')
// (9, 7, 'sp4_v_b_17')
// (9, 8, 'sp4_v_b_4')

wire n169;
// (4, 2, 'neigh_op_tnr_3')
// (4, 3, 'neigh_op_rgt_3')
// (4, 3, 'sp4_h_r_11')
// (4, 4, 'neigh_op_bnr_3')
// (5, 0, 'span12_vert_10')
// (5, 1, 'sp12_v_b_10')
// (5, 1, 'sp4_r_v_b_47')
// (5, 2, 'neigh_op_top_3')
// (5, 2, 'sp12_v_b_9')
// (5, 2, 'sp4_r_v_b_34')
// (5, 3, 'lutff_3/out')
// (5, 3, 'sp12_v_b_6')
// (5, 3, 'sp4_h_r_22')
// (5, 3, 'sp4_r_v_b_23')
// (5, 4, 'neigh_op_bot_3')
// (5, 4, 'sp12_v_b_5')
// (5, 4, 'sp4_r_v_b_10')
// (5, 5, 'sp12_v_b_2')
// (5, 5, 'sp4_r_v_b_36')
// (5, 6, 'sp12_h_r_1')
// (5, 6, 'sp12_v_b_1')
// (5, 6, 'sp4_r_v_b_25')
// (5, 7, 'sp4_r_v_b_12')
// (5, 8, 'sp4_r_v_b_1')
// (6, 0, 'span4_vert_47')
// (6, 1, 'sp4_v_b_47')
// (6, 2, 'neigh_op_tnl_3')
// (6, 2, 'sp4_v_b_34')
// (6, 3, 'neigh_op_lft_3')
// (6, 3, 'sp4_h_r_35')
// (6, 3, 'sp4_v_b_23')
// (6, 4, 'neigh_op_bnl_3')
// (6, 4, 'sp4_v_b_10')
// (6, 4, 'sp4_v_t_36')
// (6, 5, 'sp4_v_b_36')
// (6, 6, 'sp12_h_r_2')
// (6, 6, 'sp4_v_b_25')
// (6, 7, 'sp4_v_b_12')
// (6, 8, 'local_g0_1')
// (6, 8, 'lutff_6/in_1')
// (6, 8, 'sp4_h_r_1')
// (6, 8, 'sp4_v_b_1')
// (7, 3, 'sp4_h_r_46')
// (7, 4, 'sp4_r_v_b_46')
// (7, 5, 'sp4_r_v_b_35')
// (7, 6, 'sp12_h_r_5')
// (7, 6, 'sp4_r_v_b_22')
// (7, 7, 'sp4_r_v_b_11')
// (7, 8, 'sp4_h_r_12')
// (7, 8, 'sp4_r_v_b_46')
// (7, 9, 'sp4_r_v_b_35')
// (7, 10, 'sp4_r_v_b_22')
// (7, 11, 'sp4_r_v_b_11')
// (8, 3, 'sp4_h_l_46')
// (8, 3, 'sp4_v_t_46')
// (8, 4, 'sp4_v_b_46')
// (8, 5, 'sp4_v_b_35')
// (8, 6, 'local_g0_6')
// (8, 6, 'lutff_3/in_1')
// (8, 6, 'sp12_h_r_6')
// (8, 6, 'sp4_v_b_22')
// (8, 7, 'local_g0_3')
// (8, 7, 'lutff_0/in_1')
// (8, 7, 'sp4_v_b_11')
// (8, 7, 'sp4_v_t_46')
// (8, 8, 'local_g3_1')
// (8, 8, 'lutff_5/in_1')
// (8, 8, 'sp4_h_r_25')
// (8, 8, 'sp4_v_b_46')
// (8, 9, 'local_g2_3')
// (8, 9, 'lutff_6/in_1')
// (8, 9, 'sp4_v_b_35')
// (8, 10, 'sp4_v_b_22')
// (8, 11, 'sp4_v_b_11')
// (9, 5, 'sp4_r_v_b_36')
// (9, 5, 'sp4_r_v_b_42')
// (9, 6, 'local_g1_1')
// (9, 6, 'lutff_5/in_1')
// (9, 6, 'sp12_h_r_9')
// (9, 6, 'sp4_r_v_b_25')
// (9, 6, 'sp4_r_v_b_31')
// (9, 7, 'local_g3_2')
// (9, 7, 'lutff_0/in_1')
// (9, 7, 'sp4_r_v_b_12')
// (9, 7, 'sp4_r_v_b_18')
// (9, 8, 'local_g3_4')
// (9, 8, 'lutff_0/in_3')
// (9, 8, 'sp4_h_r_36')
// (9, 8, 'sp4_r_v_b_1')
// (9, 8, 'sp4_r_v_b_7')
// (9, 9, 'local_g2_4')
// (9, 9, 'lutff_5/in_1')
// (9, 9, 'sp4_r_v_b_36')
// (9, 10, 'sp4_r_v_b_25')
// (9, 11, 'sp4_r_v_b_12')
// (9, 12, 'sp4_r_v_b_1')
// (10, 4, 'sp4_v_t_36')
// (10, 4, 'sp4_v_t_42')
// (10, 5, 'sp4_v_b_36')
// (10, 5, 'sp4_v_b_42')
// (10, 6, 'sp12_h_r_10')
// (10, 6, 'sp4_v_b_25')
// (10, 6, 'sp4_v_b_31')
// (10, 7, 'sp4_v_b_12')
// (10, 7, 'sp4_v_b_18')
// (10, 8, 'sp4_h_l_36')
// (10, 8, 'sp4_v_b_1')
// (10, 8, 'sp4_v_b_7')
// (10, 8, 'sp4_v_t_36')
// (10, 9, 'sp4_v_b_36')
// (10, 10, 'sp4_v_b_25')
// (10, 11, 'sp4_v_b_12')
// (10, 12, 'sp4_v_b_1')
// (11, 6, 'sp12_h_r_13')
// (12, 6, 'sp12_h_r_14')
// (13, 6, 'span12_horz_14')

wire n170;
// (4, 3, 'lutff_1/cout')
// (4, 3, 'lutff_2/in_3')

wire n171;
// (4, 3, 'lutff_2/cout')
// (4, 3, 'lutff_3/in_3')

wire n172;
// (4, 3, 'neigh_op_tnr_5')
// (4, 4, 'neigh_op_rgt_5')
// (4, 5, 'neigh_op_bnr_5')
// (5, 1, 'sp4_r_v_b_46')
// (5, 2, 'local_g2_3')
// (5, 2, 'lutff_3/in_2')
// (5, 2, 'sp4_r_v_b_35')
// (5, 3, 'neigh_op_top_5')
// (5, 3, 'sp4_r_v_b_22')
// (5, 4, 'lutff_5/out')
// (5, 4, 'sp4_r_v_b_11')
// (5, 5, 'neigh_op_bot_5')
// (6, 0, 'span4_vert_46')
// (6, 1, 'sp4_v_b_46')
// (6, 2, 'sp4_v_b_35')
// (6, 3, 'neigh_op_tnl_5')
// (6, 3, 'sp4_v_b_22')
// (6, 4, 'neigh_op_lft_5')
// (6, 4, 'sp4_v_b_11')
// (6, 5, 'neigh_op_bnl_5')

wire n173;
// (4, 3, 'sp4_h_r_3')
// (5, 3, 'sp4_h_r_14')
// (6, 2, 'neigh_op_tnr_3')
// (6, 3, 'neigh_op_rgt_3')
// (6, 3, 'sp4_h_r_27')
// (6, 4, 'neigh_op_bnr_3')
// (7, 2, 'neigh_op_top_3')
// (7, 3, 'local_g3_6')
// (7, 3, 'lutff_1/in_2')
// (7, 3, 'lutff_3/out')
// (7, 3, 'sp4_h_r_38')
// (7, 3, 'sp4_r_v_b_39')
// (7, 4, 'local_g1_2')
// (7, 4, 'local_g1_3')
// (7, 4, 'lutff_2/in_1')
// (7, 4, 'lutff_3/in_1')
// (7, 4, 'neigh_op_bot_3')
// (7, 4, 'sp4_r_v_b_26')
// (7, 5, 'sp4_r_v_b_15')
// (7, 6, 'sp4_r_v_b_2')
// (8, 2, 'neigh_op_tnl_3')
// (8, 2, 'sp4_v_t_39')
// (8, 3, 'neigh_op_lft_3')
// (8, 3, 'sp4_h_l_38')
// (8, 3, 'sp4_v_b_39')
// (8, 4, 'neigh_op_bnl_3')
// (8, 4, 'sp4_v_b_26')
// (8, 5, 'sp4_v_b_15')
// (8, 6, 'sp4_v_b_2')

reg n174 = 0;
// (4, 4, 'neigh_op_tnr_3')
// (4, 5, 'neigh_op_rgt_3')
// (4, 6, 'neigh_op_bnr_3')
// (5, 4, 'neigh_op_top_3')
// (5, 5, 'local_g1_3')
// (5, 5, 'lutff_3/out')
// (5, 5, 'lutff_4/in_0')
// (5, 6, 'neigh_op_bot_3')
// (6, 4, 'neigh_op_tnl_3')
// (6, 5, 'neigh_op_lft_3')
// (6, 6, 'neigh_op_bnl_3')

reg n175 = 0;
// (4, 4, 'neigh_op_tnr_7')
// (4, 5, 'neigh_op_rgt_7')
// (4, 6, 'neigh_op_bnr_7')
// (5, 4, 'neigh_op_top_7')
// (5, 5, 'local_g0_7')
// (5, 5, 'lutff_2/in_1')
// (5, 5, 'lutff_7/out')
// (5, 6, 'neigh_op_bot_7')
// (6, 4, 'neigh_op_tnl_7')
// (6, 5, 'neigh_op_lft_7')
// (6, 6, 'neigh_op_bnl_7')

wire n176;
// (4, 4, 'sp12_h_r_1')
// (5, 4, 'sp12_h_r_2')
// (6, 3, 'neigh_op_tnr_7')
// (6, 4, 'neigh_op_rgt_7')
// (6, 4, 'sp12_h_r_5')
// (6, 5, 'neigh_op_bnr_7')
// (7, 3, 'neigh_op_top_7')
// (7, 4, 'lutff_7/out')
// (7, 4, 'sp12_h_r_6')
// (7, 5, 'neigh_op_bot_7')
// (8, 3, 'neigh_op_tnl_7')
// (8, 4, 'neigh_op_lft_7')
// (8, 4, 'sp12_h_r_9')
// (8, 5, 'neigh_op_bnl_7')
// (9, 4, 'local_g0_2')
// (9, 4, 'lutff_0/in_2')
// (9, 4, 'lutff_7/in_3')
// (9, 4, 'sp12_h_r_10')
// (10, 4, 'sp12_h_r_13')
// (11, 4, 'sp12_h_r_14')
// (12, 4, 'sp12_h_r_17')
// (13, 4, 'span12_horz_17')

wire n177;
// (4, 4, 'sp4_h_r_4')
// (5, 3, 'neigh_op_tnr_6')
// (5, 4, 'neigh_op_rgt_6')
// (5, 4, 'sp4_h_r_17')
// (5, 5, 'neigh_op_bnr_6')
// (6, 3, 'neigh_op_top_6')
// (6, 4, 'lutff_6/out')
// (6, 4, 'sp4_h_r_28')
// (6, 5, 'neigh_op_bot_6')
// (7, 3, 'neigh_op_tnl_6')
// (7, 4, 'local_g3_1')
// (7, 4, 'lutff_3/in_3')
// (7, 4, 'neigh_op_lft_6')
// (7, 4, 'sp4_h_r_41')
// (7, 5, 'neigh_op_bnl_6')
// (8, 4, 'sp4_h_l_41')

wire n178;
// (4, 4, 'sp4_r_v_b_42')
// (4, 5, 'sp4_r_v_b_31')
// (4, 6, 'sp4_r_v_b_18')
// (4, 7, 'sp4_r_v_b_7')
// (4, 10, 'neigh_op_tnr_1')
// (4, 11, 'neigh_op_rgt_1')
// (4, 12, 'neigh_op_bnr_1')
// (5, 0, 'span12_vert_22')
// (5, 1, 'sp12_v_b_22')
// (5, 2, 'sp12_v_b_21')
// (5, 3, 'sp12_v_b_18')
// (5, 3, 'sp4_v_t_42')
// (5, 4, 'sp12_v_b_17')
// (5, 4, 'sp4_v_b_42')
// (5, 5, 'sp12_v_b_14')
// (5, 5, 'sp4_v_b_31')
// (5, 6, 'local_g2_5')
// (5, 6, 'local_g3_5')
// (5, 6, 'lutff_0/in_2')
// (5, 6, 'lutff_3/in_3')
// (5, 6, 'lutff_4/in_3')
// (5, 6, 'lutff_5/in_1')
// (5, 6, 'lutff_7/in_2')
// (5, 6, 'sp12_v_b_13')
// (5, 6, 'sp4_v_b_18')
// (5, 7, 'local_g0_7')
// (5, 7, 'lutff_4/in_1')
// (5, 7, 'sp12_v_b_10')
// (5, 7, 'sp4_h_r_1')
// (5, 7, 'sp4_h_r_7')
// (5, 7, 'sp4_v_b_7')
// (5, 8, 'sp12_v_b_9')
// (5, 9, 'sp12_v_b_6')
// (5, 10, 'neigh_op_top_1')
// (5, 10, 'sp12_v_b_5')
// (5, 11, 'lutff_1/out')
// (5, 11, 'sp12_v_b_2')
// (5, 12, 'neigh_op_bot_1')
// (5, 12, 'sp12_v_b_1')
// (6, 7, 'local_g0_4')
// (6, 7, 'local_g1_2')
// (6, 7, 'lutff_3/in_2')
// (6, 7, 'lutff_5/in_1')
// (6, 7, 'sp4_h_r_12')
// (6, 7, 'sp4_h_r_18')
// (6, 10, 'neigh_op_tnl_1')
// (6, 11, 'neigh_op_lft_1')
// (6, 12, 'neigh_op_bnl_1')
// (7, 7, 'sp4_h_r_25')
// (7, 7, 'sp4_h_r_31')
// (8, 7, 'sp4_h_r_36')
// (8, 7, 'sp4_h_r_42')
// (9, 7, 'sp4_h_l_36')
// (9, 7, 'sp4_h_l_42')

wire n179;
// (4, 5, 'local_g0_1')
// (4, 5, 'local_g1_1')
// (4, 5, 'lutff_4/in_2')
// (4, 5, 'lutff_5/in_2')
// (4, 5, 'sp4_h_r_1')
// (5, 5, 'sp4_h_r_12')
// (6, 4, 'neigh_op_tnr_2')
// (6, 5, 'local_g3_2')
// (6, 5, 'lutff_7/in_0')
// (6, 5, 'neigh_op_rgt_2')
// (6, 5, 'sp4_h_r_25')
// (6, 6, 'neigh_op_bnr_2')
// (7, 3, 'sp4_r_v_b_45')
// (7, 4, 'neigh_op_top_2')
// (7, 4, 'sp4_r_v_b_32')
// (7, 5, 'lutff_2/out')
// (7, 5, 'sp4_h_r_36')
// (7, 5, 'sp4_r_v_b_21')
// (7, 6, 'neigh_op_bot_2')
// (7, 6, 'sp4_r_v_b_8')
// (8, 2, 'sp4_v_t_45')
// (8, 3, 'sp4_v_b_45')
// (8, 4, 'neigh_op_tnl_2')
// (8, 4, 'sp4_v_b_32')
// (8, 5, 'neigh_op_lft_2')
// (8, 5, 'sp4_h_l_36')
// (8, 5, 'sp4_v_b_21')
// (8, 6, 'neigh_op_bnl_2')
// (8, 6, 'sp4_h_r_8')
// (8, 6, 'sp4_v_b_8')
// (9, 6, 'local_g0_5')
// (9, 6, 'lutff_5/in_2')
// (9, 6, 'sp4_h_r_21')
// (10, 6, 'sp4_h_r_32')
// (11, 6, 'sp4_h_r_45')
// (12, 6, 'sp4_h_l_45')

wire n180;
// (4, 5, 'neigh_op_tnr_0')
// (4, 6, 'neigh_op_rgt_0')
// (4, 7, 'neigh_op_bnr_0')
// (5, 5, 'neigh_op_top_0')
// (5, 6, 'local_g1_0')
// (5, 6, 'lutff_0/out')
// (5, 6, 'lutff_5/in_2')
// (5, 6, 'lutff_6/in_3')
// (5, 7, 'local_g0_0')
// (5, 7, 'local_g1_0')
// (5, 7, 'lutff_1/in_1')
// (5, 7, 'lutff_6/in_3')
// (5, 7, 'neigh_op_bot_0')
// (6, 5, 'neigh_op_tnl_0')
// (6, 6, 'neigh_op_lft_0')
// (6, 7, 'neigh_op_bnl_0')

wire n181;
// (4, 5, 'neigh_op_tnr_1')
// (4, 6, 'local_g2_1')
// (4, 6, 'lutff_2/in_3')
// (4, 6, 'neigh_op_rgt_1')
// (4, 7, 'neigh_op_bnr_1')
// (5, 5, 'neigh_op_top_1')
// (5, 6, 'lutff_1/out')
// (5, 7, 'neigh_op_bot_1')
// (6, 5, 'neigh_op_tnl_1')
// (6, 6, 'neigh_op_lft_1')
// (6, 7, 'neigh_op_bnl_1')

wire n182;
// (4, 5, 'neigh_op_tnr_2')
// (4, 6, 'local_g3_2')
// (4, 6, 'lutff_0/in_3')
// (4, 6, 'neigh_op_rgt_2')
// (4, 7, 'neigh_op_bnr_2')
// (5, 5, 'neigh_op_top_2')
// (5, 6, 'lutff_2/out')
// (5, 7, 'neigh_op_bot_2')
// (6, 5, 'neigh_op_tnl_2')
// (6, 6, 'neigh_op_lft_2')
// (6, 7, 'neigh_op_bnl_2')

wire n183;
// (4, 5, 'neigh_op_tnr_4')
// (4, 6, 'local_g2_4')
// (4, 6, 'lutff_3/in_1')
// (4, 6, 'neigh_op_rgt_4')
// (4, 7, 'neigh_op_bnr_4')
// (5, 5, 'neigh_op_top_4')
// (5, 6, 'lutff_4/out')
// (5, 7, 'neigh_op_bot_4')
// (6, 5, 'neigh_op_tnl_4')
// (6, 6, 'neigh_op_lft_4')
// (6, 7, 'neigh_op_bnl_4')

wire n184;
// (4, 5, 'neigh_op_tnr_7')
// (4, 6, 'local_g3_7')
// (4, 6, 'lutff_0/in_0')
// (4, 6, 'lutff_6/in_2')
// (4, 6, 'neigh_op_rgt_7')
// (4, 7, 'local_g0_7')
// (4, 7, 'local_g1_7')
// (4, 7, 'lutff_0/in_3')
// (4, 7, 'lutff_5/in_3')
// (4, 7, 'neigh_op_bnr_7')
// (5, 5, 'neigh_op_top_7')
// (5, 6, 'local_g1_7')
// (5, 6, 'lutff_4/in_2')
// (5, 6, 'lutff_7/out')
// (5, 7, 'neigh_op_bot_7')
// (6, 5, 'neigh_op_tnl_7')
// (6, 6, 'neigh_op_lft_7')
// (6, 7, 'neigh_op_bnl_7')

wire n185;
// (4, 5, 'sp4_r_v_b_42')
// (4, 6, 'neigh_op_tnr_1')
// (4, 6, 'sp4_r_v_b_31')
// (4, 7, 'neigh_op_rgt_1')
// (4, 7, 'sp4_r_v_b_18')
// (4, 8, 'local_g1_1')
// (4, 8, 'lutff_2/in_2')
// (4, 8, 'lutff_6/in_0')
// (4, 8, 'neigh_op_bnr_1')
// (4, 8, 'sp4_r_v_b_7')
// (5, 0, 'span12_vert_14')
// (5, 1, 'sp12_v_b_14')
// (5, 2, 'sp12_v_b_13')
// (5, 3, 'sp12_v_b_10')
// (5, 4, 'sp12_v_b_9')
// (5, 4, 'sp4_v_t_42')
// (5, 5, 'sp12_v_b_6')
// (5, 5, 'sp4_v_b_42')
// (5, 6, 'neigh_op_top_1')
// (5, 6, 'sp12_v_b_5')
// (5, 6, 'sp4_v_b_31')
// (5, 7, 'lutff_1/out')
// (5, 7, 'sp12_v_b_2')
// (5, 7, 'sp4_v_b_18')
// (5, 8, 'local_g0_7')
// (5, 8, 'local_g3_1')
// (5, 8, 'lutff_4/in_2')
// (5, 8, 'lutff_5/in_0')
// (5, 8, 'neigh_op_bot_1')
// (5, 8, 'sp12_v_b_1')
// (5, 8, 'sp4_v_b_7')
// (6, 6, 'neigh_op_tnl_1')
// (6, 7, 'neigh_op_lft_1')
// (6, 8, 'neigh_op_bnl_1')

wire n186;
// (4, 6, 'local_g2_0')
// (4, 6, 'local_g3_0')
// (4, 6, 'lutff_0/in_1')
// (4, 6, 'lutff_6/in_0')
// (4, 6, 'neigh_op_tnr_0')
// (4, 7, 'local_g2_0')
// (4, 7, 'local_g3_0')
// (4, 7, 'lutff_1/in_3')
// (4, 7, 'lutff_2/in_3')
// (4, 7, 'neigh_op_rgt_0')
// (4, 8, 'neigh_op_bnr_0')
// (5, 6, 'local_g0_0')
// (5, 6, 'lutff_4/in_0')
// (5, 6, 'neigh_op_top_0')
// (5, 7, 'lutff_0/out')
// (5, 8, 'neigh_op_bot_0')
// (6, 6, 'neigh_op_tnl_0')
// (6, 7, 'neigh_op_lft_0')
// (6, 8, 'neigh_op_bnl_0')

wire n187;
// (4, 6, 'neigh_op_tnr_3')
// (4, 7, 'neigh_op_rgt_3')
// (4, 8, 'neigh_op_bnr_3')
// (5, 6, 'neigh_op_top_3')
// (5, 7, 'local_g1_3')
// (5, 7, 'lutff_3/out')
// (5, 7, 'lutff_4/in_0')
// (5, 7, 'lutff_6/in_0')
// (5, 8, 'neigh_op_bot_3')
// (6, 6, 'neigh_op_tnl_3')
// (6, 7, 'neigh_op_lft_3')
// (6, 8, 'neigh_op_bnl_3')

wire n188;
// (4, 6, 'neigh_op_tnr_4')
// (4, 7, 'neigh_op_rgt_4')
// (4, 8, 'local_g1_4')
// (4, 8, 'lutff_4/in_3')
// (4, 8, 'lutff_5/in_2')
// (4, 8, 'neigh_op_bnr_4')
// (5, 6, 'neigh_op_top_4')
// (5, 6, 'sp4_r_v_b_36')
// (5, 7, 'lutff_4/out')
// (5, 7, 'sp4_r_v_b_25')
// (5, 8, 'neigh_op_bot_4')
// (5, 8, 'sp4_r_v_b_12')
// (5, 9, 'local_g1_1')
// (5, 9, 'lutff_5/in_3')
// (5, 9, 'sp4_r_v_b_1')
// (6, 5, 'sp4_v_t_36')
// (6, 6, 'neigh_op_tnl_4')
// (6, 6, 'sp4_v_b_36')
// (6, 7, 'neigh_op_lft_4')
// (6, 7, 'sp4_v_b_25')
// (6, 8, 'neigh_op_bnl_4')
// (6, 8, 'sp4_v_b_12')
// (6, 9, 'sp4_v_b_1')

wire n189;
// (4, 6, 'neigh_op_tnr_5')
// (4, 7, 'neigh_op_rgt_5')
// (4, 8, 'neigh_op_bnr_5')
// (5, 6, 'local_g0_5')
// (5, 6, 'local_g1_5')
// (5, 6, 'lutff_1/in_3')
// (5, 6, 'lutff_2/in_1')
// (5, 6, 'neigh_op_top_5')
// (5, 7, 'lutff_5/out')
// (5, 8, 'local_g0_5')
// (5, 8, 'local_g1_5')
// (5, 8, 'lutff_2/in_1')
// (5, 8, 'lutff_3/in_3')
// (5, 8, 'neigh_op_bot_5')
// (6, 6, 'neigh_op_tnl_5')
// (6, 7, 'neigh_op_lft_5')
// (6, 8, 'neigh_op_bnl_5')

wire n190;
// (4, 6, 'neigh_op_tnr_6')
// (4, 7, 'neigh_op_rgt_6')
// (4, 8, 'local_g0_6')
// (4, 8, 'local_g1_6')
// (4, 8, 'lutff_5/in_3')
// (4, 8, 'lutff_6/in_3')
// (4, 8, 'neigh_op_bnr_6')
// (5, 6, 'neigh_op_top_6')
// (5, 7, 'lutff_6/out')
// (5, 8, 'neigh_op_bot_6')
// (6, 6, 'neigh_op_tnl_6')
// (6, 7, 'neigh_op_lft_6')
// (6, 8, 'neigh_op_bnl_6')

wire n191;
// (4, 6, 'neigh_op_tnr_7')
// (4, 7, 'neigh_op_rgt_7')
// (4, 8, 'neigh_op_bnr_7')
// (5, 6, 'neigh_op_top_7')
// (5, 7, 'lutff_7/out')
// (5, 8, 'local_g1_7')
// (5, 8, 'lutff_2/in_0')
// (5, 8, 'lutff_6/in_0')
// (5, 8, 'neigh_op_bot_7')
// (6, 6, 'neigh_op_tnl_7')
// (6, 7, 'neigh_op_lft_7')
// (6, 8, 'neigh_op_bnl_7')

wire n192;
// (4, 7, 'neigh_op_tnr_0')
// (4, 8, 'neigh_op_rgt_0')
// (4, 9, 'neigh_op_bnr_0')
// (5, 7, 'neigh_op_top_0')
// (5, 8, 'local_g2_0')
// (5, 8, 'lutff_0/out')
// (5, 8, 'lutff_5/in_3')
// (5, 9, 'neigh_op_bot_0')
// (6, 7, 'neigh_op_tnl_0')
// (6, 8, 'neigh_op_lft_0')
// (6, 9, 'neigh_op_bnl_0')

wire n193;
// (4, 7, 'neigh_op_tnr_1')
// (4, 8, 'neigh_op_rgt_1')
// (4, 9, 'neigh_op_bnr_1')
// (5, 7, 'neigh_op_top_1')
// (5, 8, 'local_g2_1')
// (5, 8, 'lutff_0/in_1')
// (5, 8, 'lutff_1/out')
// (5, 8, 'lutff_6/in_3')
// (5, 9, 'neigh_op_bot_1')
// (6, 7, 'neigh_op_tnl_1')
// (6, 8, 'neigh_op_lft_1')
// (6, 9, 'neigh_op_bnl_1')

wire n194;
// (4, 7, 'neigh_op_tnr_2')
// (4, 8, 'local_g2_2')
// (4, 8, 'local_g3_2')
// (4, 8, 'lutff_0/in_3')
// (4, 8, 'lutff_4/in_2')
// (4, 8, 'neigh_op_rgt_2')
// (4, 9, 'neigh_op_bnr_2')
// (5, 7, 'neigh_op_top_2')
// (5, 8, 'lutff_2/out')
// (5, 9, 'neigh_op_bot_2')
// (6, 7, 'neigh_op_tnl_2')
// (6, 8, 'neigh_op_lft_2')
// (6, 9, 'neigh_op_bnl_2')

wire n195;
// (4, 7, 'neigh_op_tnr_3')
// (4, 8, 'local_g2_3')
// (4, 8, 'lutff_2/in_3')
// (4, 8, 'lutff_3/in_2')
// (4, 8, 'lutff_6/in_1')
// (4, 8, 'neigh_op_rgt_3')
// (4, 9, 'neigh_op_bnr_3')
// (5, 7, 'neigh_op_top_3')
// (5, 8, 'local_g0_3')
// (5, 8, 'lutff_3/out')
// (5, 8, 'lutff_4/in_3')
// (5, 9, 'neigh_op_bot_3')
// (6, 7, 'neigh_op_tnl_3')
// (6, 8, 'neigh_op_lft_3')
// (6, 9, 'neigh_op_bnl_3')

wire n196;
// (4, 7, 'neigh_op_tnr_4')
// (4, 8, 'neigh_op_rgt_4')
// (4, 9, 'neigh_op_bnr_4')
// (5, 7, 'neigh_op_top_4')
// (5, 7, 'sp4_r_v_b_36')
// (5, 8, 'lutff_4/out')
// (5, 8, 'sp4_r_v_b_25')
// (5, 9, 'neigh_op_bot_4')
// (5, 9, 'sp4_r_v_b_12')
// (5, 10, 'sp4_r_v_b_1')
// (6, 6, 'sp4_v_t_36')
// (6, 7, 'neigh_op_tnl_4')
// (6, 7, 'sp4_v_b_36')
// (6, 8, 'neigh_op_lft_4')
// (6, 8, 'sp4_v_b_25')
// (6, 9, 'neigh_op_bnl_4')
// (6, 9, 'sp4_v_b_12')
// (6, 10, 'local_g0_7')
// (6, 10, 'local_g1_1')
// (6, 10, 'lutff_1/in_3')
// (6, 10, 'lutff_4/in_3')
// (6, 10, 'sp4_h_r_7')
// (6, 10, 'sp4_v_b_1')
// (7, 10, 'local_g1_2')
// (7, 10, 'lutff_1/in_2')
// (7, 10, 'sp4_h_r_18')
// (8, 10, 'sp4_h_r_31')
// (9, 10, 'sp4_h_r_42')
// (10, 10, 'sp4_h_l_42')
// (10, 10, 'sp4_h_r_10')
// (11, 10, 'local_g0_7')
// (11, 10, 'lutff_2/in_3')
// (11, 10, 'sp4_h_r_23')
// (12, 10, 'sp4_h_r_34')
// (13, 10, 'span4_horz_34')

wire n197;
// (4, 7, 'neigh_op_tnr_5')
// (4, 8, 'neigh_op_rgt_5')
// (4, 8, 'sp4_r_v_b_42')
// (4, 9, 'local_g1_7')
// (4, 9, 'lutff_3/in_3')
// (4, 9, 'neigh_op_bnr_5')
// (4, 9, 'sp4_r_v_b_31')
// (4, 9, 'sp4_r_v_b_41')
// (4, 10, 'local_g0_4')
// (4, 10, 'local_g3_2')
// (4, 10, 'lutff_0/in_2')
// (4, 10, 'lutff_3/in_3')
// (4, 10, 'lutff_4/in_3')
// (4, 10, 'sp4_r_v_b_18')
// (4, 10, 'sp4_r_v_b_28')
// (4, 11, 'sp4_r_v_b_17')
// (4, 11, 'sp4_r_v_b_7')
// (4, 12, 'sp4_r_v_b_4')
// (5, 5, 'sp4_r_v_b_46')
// (5, 6, 'sp4_r_v_b_35')
// (5, 7, 'neigh_op_top_5')
// (5, 7, 'sp4_r_v_b_22')
// (5, 7, 'sp4_v_t_42')
// (5, 8, 'lutff_5/out')
// (5, 8, 'sp4_h_r_10')
// (5, 8, 'sp4_r_v_b_11')
// (5, 8, 'sp4_v_b_42')
// (5, 8, 'sp4_v_t_41')
// (5, 9, 'neigh_op_bot_5')
// (5, 9, 'sp4_v_b_31')
// (5, 9, 'sp4_v_b_41')
// (5, 10, 'sp4_v_b_18')
// (5, 10, 'sp4_v_b_28')
// (5, 11, 'sp4_v_b_17')
// (5, 11, 'sp4_v_b_7')
// (5, 12, 'sp4_v_b_4')
// (6, 4, 'sp4_v_t_46')
// (6, 5, 'sp4_v_b_46')
// (6, 6, 'local_g2_3')
// (6, 6, 'lutff_6/in_3')
// (6, 6, 'sp4_v_b_35')
// (6, 7, 'neigh_op_tnl_5')
// (6, 7, 'sp4_v_b_22')
// (6, 8, 'local_g0_5')
// (6, 8, 'lutff_0/in_1')
// (6, 8, 'lutff_3/in_2')
// (6, 8, 'neigh_op_lft_5')
// (6, 8, 'sp4_h_r_23')
// (6, 8, 'sp4_v_b_11')
// (6, 9, 'neigh_op_bnl_5')
// (7, 8, 'sp4_h_r_34')
// (8, 8, 'sp4_h_r_47')
// (9, 8, 'sp4_h_l_47')

wire n198;
// (4, 7, 'neigh_op_tnr_6')
// (4, 8, 'local_g2_6')
// (4, 8, 'lutff_7/in_3')
// (4, 8, 'neigh_op_rgt_6')
// (4, 9, 'neigh_op_bnr_6')
// (5, 7, 'neigh_op_top_6')
// (5, 8, 'local_g3_6')
// (5, 8, 'lutff_4/in_1')
// (5, 8, 'lutff_6/out')
// (5, 9, 'neigh_op_bot_6')
// (6, 7, 'neigh_op_tnl_6')
// (6, 8, 'neigh_op_lft_6')
// (6, 9, 'neigh_op_bnl_6')

reg n199 = 0;
// (4, 7, 'neigh_op_tnr_7')
// (4, 8, 'neigh_op_rgt_7')
// (4, 8, 'sp4_h_r_3')
// (4, 9, 'neigh_op_bnr_7')
// (5, 7, 'neigh_op_top_7')
// (5, 8, 'lutff_7/out')
// (5, 8, 'sp4_h_r_14')
// (5, 9, 'neigh_op_bot_7')
// (6, 7, 'neigh_op_tnl_7')
// (6, 8, 'neigh_op_lft_7')
// (6, 8, 'sp4_h_r_27')
// (6, 9, 'neigh_op_bnl_7')
// (7, 8, 'local_g2_6')
// (7, 8, 'lutff_7/in_1')
// (7, 8, 'sp4_h_r_38')
// (8, 8, 'sp4_h_l_38')

wire n200;
// (4, 7, 'sp4_h_r_8')
// (5, 6, 'neigh_op_tnr_0')
// (5, 6, 'sp4_r_v_b_45')
// (5, 7, 'local_g0_3')
// (5, 7, 'local_g1_5')
// (5, 7, 'lutff_1/in_2')
// (5, 7, 'lutff_4/in_2')
// (5, 7, 'lutff_6/in_2')
// (5, 7, 'neigh_op_rgt_0')
// (5, 7, 'sp4_h_r_21')
// (5, 7, 'sp4_r_v_b_32')
// (5, 8, 'neigh_op_bnr_0')
// (5, 8, 'sp4_r_v_b_21')
// (5, 9, 'sp4_r_v_b_8')
// (6, 5, 'sp4_v_t_45')
// (6, 6, 'neigh_op_top_0')
// (6, 6, 'sp4_v_b_45')
// (6, 7, 'local_g2_0')
// (6, 7, 'lutff_0/out')
// (6, 7, 'lutff_3/in_3')
// (6, 7, 'sp4_h_r_32')
// (6, 7, 'sp4_v_b_32')
// (6, 8, 'neigh_op_bot_0')
// (6, 8, 'sp4_v_b_21')
// (6, 9, 'sp4_v_b_8')
// (7, 6, 'neigh_op_tnl_0')
// (7, 7, 'neigh_op_lft_0')
// (7, 7, 'sp4_h_r_45')
// (7, 8, 'neigh_op_bnl_0')
// (8, 7, 'sp4_h_l_45')

wire n201;
// (4, 8, 'neigh_op_tnr_0')
// (4, 9, 'neigh_op_rgt_0')
// (4, 10, 'neigh_op_bnr_0')
// (5, 0, 'span12_vert_16')
// (5, 1, 'sp12_v_b_16')
// (5, 2, 'sp12_v_b_15')
// (5, 3, 'sp12_v_b_12')
// (5, 3, 'sp4_r_v_b_41')
// (5, 4, 'sp12_v_b_11')
// (5, 4, 'sp4_r_v_b_28')
// (5, 5, 'sp12_v_b_8')
// (5, 5, 'sp4_r_v_b_17')
// (5, 6, 'local_g1_4')
// (5, 6, 'local_g3_7')
// (5, 6, 'lutff_0/in_1')
// (5, 6, 'lutff_1/in_2')
// (5, 6, 'lutff_2/in_0')
// (5, 6, 'lutff_3/in_2')
// (5, 6, 'lutff_7/in_1')
// (5, 6, 'sp12_v_b_7')
// (5, 6, 'sp4_r_v_b_4')
// (5, 7, 'local_g3_1')
// (5, 7, 'lutff_0/in_2')
// (5, 7, 'sp12_v_b_4')
// (5, 7, 'sp4_r_v_b_37')
// (5, 7, 'sp4_r_v_b_41')
// (5, 8, 'local_g1_4')
// (5, 8, 'lutff_0/in_3')
// (5, 8, 'lutff_6/in_1')
// (5, 8, 'neigh_op_top_0')
// (5, 8, 'sp12_v_b_3')
// (5, 8, 'sp4_r_v_b_24')
// (5, 8, 'sp4_r_v_b_28')
// (5, 9, 'lutff_0/out')
// (5, 9, 'sp12_v_b_0')
// (5, 9, 'sp4_r_v_b_13')
// (5, 9, 'sp4_r_v_b_17')
// (5, 10, 'neigh_op_bot_0')
// (5, 10, 'sp4_r_v_b_0')
// (5, 10, 'sp4_r_v_b_4')
// (6, 2, 'sp4_v_t_41')
// (6, 3, 'sp4_v_b_41')
// (6, 4, 'sp4_v_b_28')
// (6, 5, 'sp4_v_b_17')
// (6, 6, 'sp4_v_b_4')
// (6, 6, 'sp4_v_t_37')
// (6, 6, 'sp4_v_t_41')
// (6, 7, 'local_g2_5')
// (6, 7, 'lutff_2/in_1')
// (6, 7, 'sp4_v_b_37')
// (6, 7, 'sp4_v_b_41')
// (6, 8, 'neigh_op_tnl_0')
// (6, 8, 'sp4_v_b_24')
// (6, 8, 'sp4_v_b_28')
// (6, 9, 'neigh_op_lft_0')
// (6, 9, 'sp4_v_b_13')
// (6, 9, 'sp4_v_b_17')
// (6, 10, 'neigh_op_bnl_0')
// (6, 10, 'sp4_v_b_0')
// (6, 10, 'sp4_v_b_4')

wire n202;
// (4, 8, 'neigh_op_tnr_2')
// (4, 9, 'neigh_op_rgt_2')
// (4, 9, 'sp4_h_r_9')
// (4, 9, 'sp4_r_v_b_36')
// (4, 10, 'neigh_op_bnr_2')
// (4, 10, 'sp4_r_v_b_25')
// (4, 11, 'sp4_r_v_b_12')
// (4, 12, 'sp4_r_v_b_1')
// (4, 13, 'sp4_h_r_2')
// (5, 0, 'span12_vert_20')
// (5, 1, 'sp12_v_b_20')
// (5, 2, 'sp12_v_b_19')
// (5, 3, 'sp12_v_b_16')
// (5, 4, 'sp12_v_b_15')
// (5, 5, 'sp12_v_b_12')
// (5, 6, 'sp12_v_b_11')
// (5, 7, 'sp12_v_b_8')
// (5, 8, 'neigh_op_top_2')
// (5, 8, 'sp12_v_b_7')
// (5, 8, 'sp4_v_t_36')
// (5, 9, 'lutff_2/out')
// (5, 9, 'sp12_v_b_4')
// (5, 9, 'sp4_h_r_20')
// (5, 9, 'sp4_v_b_36')
// (5, 10, 'neigh_op_bot_2')
// (5, 10, 'sp12_v_b_3')
// (5, 10, 'sp4_v_b_25')
// (5, 11, 'local_g2_0')
// (5, 11, 'lutff_2/in_0')
// (5, 11, 'sp12_h_r_0')
// (5, 11, 'sp12_v_b_0')
// (5, 11, 'sp4_v_b_12')
// (5, 12, 'local_g0_7')
// (5, 12, 'local_g1_1')
// (5, 12, 'lutff_0/in_0')
// (5, 12, 'lutff_6/in_3')
// (5, 12, 'lutff_7/in_3')
// (5, 12, 'sp4_h_r_7')
// (5, 12, 'sp4_v_b_1')
// (5, 13, 'sp4_h_r_15')
// (6, 8, 'neigh_op_tnl_2')
// (6, 9, 'neigh_op_lft_2')
// (6, 9, 'sp4_h_r_33')
// (6, 10, 'neigh_op_bnl_2')
// (6, 11, 'local_g0_3')
// (6, 11, 'lutff_1/in_0')
// (6, 11, 'sp12_h_r_3')
// (6, 12, 'local_g0_2')
// (6, 12, 'lutff_7/in_3')
// (6, 12, 'sp4_h_r_18')
// (6, 13, 'local_g2_2')
// (6, 13, 'lutff_0/in_0')
// (6, 13, 'lutff_3/in_3')
// (6, 13, 'sp4_h_r_26')
// (7, 6, 'sp4_r_v_b_44')
// (7, 7, 'sp4_r_v_b_33')
// (7, 8, 'sp4_r_v_b_20')
// (7, 9, 'local_g2_1')
// (7, 9, 'local_g2_4')
// (7, 9, 'lutff_0/in_3')
// (7, 9, 'lutff_1/in_0')
// (7, 9, 'lutff_6/in_3')
// (7, 9, 'lutff_7/in_3')
// (7, 9, 'sp4_h_r_44')
// (7, 9, 'sp4_r_v_b_9')
// (7, 10, 'sp4_r_v_b_39')
// (7, 11, 'sp12_h_r_4')
// (7, 11, 'sp4_r_v_b_26')
// (7, 12, 'local_g3_7')
// (7, 12, 'lutff_0/in_0')
// (7, 12, 'lutff_5/in_3')
// (7, 12, 'sp4_h_r_31')
// (7, 12, 'sp4_r_v_b_15')
// (7, 13, 'local_g1_2')
// (7, 13, 'local_g3_7')
// (7, 13, 'lutff_1/in_0')
// (7, 13, 'lutff_7/in_3')
// (7, 13, 'sp4_h_r_39')
// (7, 13, 'sp4_r_v_b_2')
// (8, 5, 'sp4_v_t_44')
// (8, 6, 'sp4_v_b_44')
// (8, 7, 'sp4_v_b_33')
// (8, 8, 'sp4_v_b_20')
// (8, 9, 'sp4_h_l_44')
// (8, 9, 'sp4_v_b_9')
// (8, 9, 'sp4_v_t_39')
// (8, 10, 'sp4_v_b_39')
// (8, 11, 'sp12_h_r_7')
// (8, 11, 'sp4_v_b_26')
// (8, 12, 'sp4_h_r_42')
// (8, 12, 'sp4_v_b_15')
// (8, 13, 'sp4_h_l_39')
// (8, 13, 'sp4_v_b_2')
// (9, 11, 'sp12_h_r_8')
// (9, 12, 'sp4_h_l_42')
// (10, 11, 'sp12_h_r_11')
// (11, 11, 'sp12_h_r_12')
// (12, 11, 'sp12_h_r_15')
// (13, 11, 'span12_horz_15')

wire n203;
// (4, 8, 'neigh_op_tnr_4')
// (4, 9, 'neigh_op_rgt_4')
// (4, 10, 'neigh_op_bnr_4')
// (5, 6, 'sp4_r_v_b_44')
// (5, 7, 'local_g0_2')
// (5, 7, 'lutff_2/in_2')
// (5, 7, 'lutff_5/in_3')
// (5, 7, 'sp4_r_v_b_33')
// (5, 8, 'neigh_op_top_4')
// (5, 8, 'sp4_r_v_b_20')
// (5, 9, 'lutff_4/out')
// (5, 9, 'sp4_r_v_b_9')
// (5, 10, 'neigh_op_bot_4')
// (6, 5, 'sp4_v_t_44')
// (6, 6, 'sp4_v_b_44')
// (6, 7, 'sp4_v_b_33')
// (6, 8, 'neigh_op_tnl_4')
// (6, 8, 'sp4_v_b_20')
// (6, 9, 'neigh_op_lft_4')
// (6, 9, 'sp4_v_b_9')
// (6, 10, 'neigh_op_bnl_4')

wire n204;
// (4, 8, 'neigh_op_tnr_5')
// (4, 9, 'neigh_op_rgt_5')
// (4, 10, 'neigh_op_bnr_5')
// (5, 8, 'neigh_op_top_5')
// (5, 9, 'lutff_5/out')
// (5, 10, 'neigh_op_bot_5')
// (6, 8, 'neigh_op_tnl_5')
// (6, 9, 'local_g0_5')
// (6, 9, 'lutff_2/in_3')
// (6, 9, 'neigh_op_lft_5')
// (6, 10, 'neigh_op_bnl_5')

wire n205;
// (4, 8, 'neigh_op_tnr_6')
// (4, 9, 'neigh_op_rgt_6')
// (4, 10, 'neigh_op_bnr_6')
// (5, 3, 'sp12_v_t_23')
// (5, 4, 'sp12_v_b_23')
// (5, 5, 'sp12_v_b_20')
// (5, 6, 'local_g2_3')
// (5, 6, 'lutff_1/in_0')
// (5, 6, 'lutff_2/in_3')
// (5, 6, 'lutff_7/in_0')
// (5, 6, 'sp12_v_b_19')
// (5, 7, 'local_g3_0')
// (5, 7, 'lutff_0/in_1')
// (5, 7, 'sp12_v_b_16')
// (5, 8, 'local_g1_6')
// (5, 8, 'lutff_1/in_2')
// (5, 8, 'lutff_2/in_3')
// (5, 8, 'lutff_3/in_0')
// (5, 8, 'neigh_op_top_6')
// (5, 8, 'sp12_v_b_15')
// (5, 9, 'lutff_6/out')
// (5, 9, 'sp12_v_b_12')
// (5, 10, 'neigh_op_bot_6')
// (5, 10, 'sp12_v_b_11')
// (5, 11, 'sp12_v_b_8')
// (5, 12, 'sp12_v_b_7')
// (5, 13, 'sp12_v_b_4')
// (5, 14, 'sp12_v_b_3')
// (5, 15, 'sp12_v_b_0')
// (6, 8, 'neigh_op_tnl_6')
// (6, 9, 'neigh_op_lft_6')
// (6, 10, 'neigh_op_bnl_6')

reg n206 = 0;
// (4, 9, 'neigh_op_tnr_1')
// (4, 10, 'neigh_op_rgt_1')
// (4, 11, 'local_g0_1')
// (4, 11, 'lutff_2/in_1')
// (4, 11, 'neigh_op_bnr_1')
// (5, 9, 'neigh_op_top_1')
// (5, 10, 'lutff_1/out')
// (5, 11, 'neigh_op_bot_1')
// (6, 9, 'neigh_op_tnl_1')
// (6, 10, 'neigh_op_lft_1')
// (6, 11, 'neigh_op_bnl_1')

reg n207 = 0;
// (4, 9, 'neigh_op_tnr_6')
// (4, 10, 'neigh_op_rgt_6')
// (4, 11, 'neigh_op_bnr_6')
// (5, 8, 'sp4_r_v_b_37')
// (5, 9, 'neigh_op_top_6')
// (5, 9, 'sp4_r_v_b_24')
// (5, 10, 'lutff_6/out')
// (5, 10, 'sp4_r_v_b_13')
// (5, 11, 'neigh_op_bot_6')
// (5, 11, 'sp4_r_v_b_0')
// (6, 7, 'sp4_v_t_37')
// (6, 8, 'sp4_v_b_37')
// (6, 9, 'neigh_op_tnl_6')
// (6, 9, 'sp4_v_b_24')
// (6, 10, 'local_g1_5')
// (6, 10, 'lutff_3/in_1')
// (6, 10, 'neigh_op_lft_6')
// (6, 10, 'sp4_v_b_13')
// (6, 11, 'neigh_op_bnl_6')
// (6, 11, 'sp4_v_b_0')

reg n208 = 0;
// (4, 9, 'neigh_op_tnr_7')
// (4, 10, 'neigh_op_rgt_7')
// (4, 11, 'neigh_op_bnr_7')
// (5, 9, 'neigh_op_top_7')
// (5, 10, 'lutff_7/out')
// (5, 11, 'neigh_op_bot_7')
// (6, 9, 'neigh_op_tnl_7')
// (6, 10, 'neigh_op_lft_7')
// (6, 11, 'local_g3_7')
// (6, 11, 'lutff_3/in_1')
// (6, 11, 'neigh_op_bnl_7')

reg n209 = 0;
// (4, 9, 'sp12_h_r_1')
// (5, 9, 'sp12_h_r_2')
// (6, 9, 'sp12_h_r_5')
// (7, 9, 'sp12_h_r_6')
// (8, 8, 'neigh_op_tnr_1')
// (8, 9, 'neigh_op_rgt_1')
// (8, 9, 'sp12_h_r_9')
// (8, 10, 'neigh_op_bnr_1')
// (9, 8, 'neigh_op_top_1')
// (9, 9, 'lutff_1/out')
// (9, 9, 'sp12_h_r_10')
// (9, 10, 'neigh_op_bot_1')
// (10, 8, 'neigh_op_tnl_1')
// (10, 9, 'neigh_op_lft_1')
// (10, 9, 'sp12_h_r_13')
// (10, 10, 'neigh_op_bnl_1')
// (11, 9, 'local_g1_6')
// (11, 9, 'lutff_7/in_0')
// (11, 9, 'sp12_h_r_14')
// (12, 9, 'sp12_h_r_17')
// (13, 9, 'span12_horz_17')

wire n210;
// (4, 9, 'sp4_r_v_b_39')
// (4, 10, 'sp4_r_v_b_26')
// (4, 11, 'neigh_op_tnr_1')
// (4, 11, 'sp4_r_v_b_15')
// (4, 12, 'neigh_op_rgt_1')
// (4, 12, 'sp4_r_v_b_2')
// (4, 13, 'neigh_op_bnr_1')
// (5, 8, 'sp4_v_t_39')
// (5, 9, 'sp4_v_b_39')
// (5, 10, 'sp4_v_b_26')
// (5, 11, 'local_g0_7')
// (5, 11, 'lutff_2/in_3')
// (5, 11, 'neigh_op_top_1')
// (5, 11, 'sp4_v_b_15')
// (5, 12, 'lutff_1/out')
// (5, 12, 'sp4_v_b_2')
// (5, 13, 'neigh_op_bot_1')
// (6, 11, 'neigh_op_tnl_1')
// (6, 12, 'neigh_op_lft_1')
// (6, 13, 'neigh_op_bnl_1')

wire n211;
// (4, 9, 'sp4_r_v_b_45')
// (4, 10, 'sp4_r_v_b_32')
// (4, 11, 'sp4_r_v_b_21')
// (4, 12, 'sp4_r_v_b_8')
// (5, 8, 'sp4_v_t_45')
// (5, 9, 'sp4_v_b_45')
// (5, 10, 'sp4_v_b_32')
// (5, 11, 'local_g1_5')
// (5, 11, 'lutff_1/in_3')
// (5, 11, 'sp4_v_b_21')
// (5, 12, 'sp4_h_r_8')
// (5, 12, 'sp4_v_b_8')
// (6, 11, 'neigh_op_tnr_0')
// (6, 12, 'neigh_op_rgt_0')
// (6, 12, 'sp4_h_r_21')
// (6, 13, 'neigh_op_bnr_0')
// (7, 11, 'neigh_op_top_0')
// (7, 12, 'lutff_0/out')
// (7, 12, 'sp4_h_r_32')
// (7, 13, 'neigh_op_bot_0')
// (8, 11, 'neigh_op_tnl_0')
// (8, 12, 'neigh_op_lft_0')
// (8, 12, 'sp4_h_r_45')
// (8, 13, 'neigh_op_bnl_0')
// (9, 12, 'sp4_h_l_45')

wire n212;
// (4, 10, 'neigh_op_tnr_2')
// (4, 11, 'neigh_op_rgt_2')
// (4, 12, 'neigh_op_bnr_2')
// (5, 1, 'sp12_v_t_23')
// (5, 2, 'sp12_v_b_23')
// (5, 3, 'sp12_v_b_20')
// (5, 4, 'sp12_v_b_19')
// (5, 5, 'sp12_v_b_16')
// (5, 6, 'sp12_v_b_15')
// (5, 7, 'sp12_v_b_12')
// (5, 8, 'sp12_v_b_11')
// (5, 8, 'sp4_r_v_b_40')
// (5, 9, 'local_g1_5')
// (5, 9, 'local_g3_0')
// (5, 9, 'lutff_0/in_0')
// (5, 9, 'lutff_6/in_1')
// (5, 9, 'sp12_v_b_8')
// (5, 9, 'sp4_r_v_b_29')
// (5, 10, 'neigh_op_top_2')
// (5, 10, 'sp12_v_b_7')
// (5, 10, 'sp4_r_v_b_16')
// (5, 11, 'local_g1_2')
// (5, 11, 'lutff_1/in_0')
// (5, 11, 'lutff_2/out')
// (5, 11, 'sp12_v_b_4')
// (5, 11, 'sp4_r_v_b_5')
// (5, 12, 'neigh_op_bot_2')
// (5, 12, 'sp12_v_b_3')
// (5, 13, 'sp12_v_b_0')
// (6, 7, 'sp4_v_t_40')
// (6, 8, 'sp4_v_b_40')
// (6, 9, 'sp4_v_b_29')
// (6, 10, 'neigh_op_tnl_2')
// (6, 10, 'sp4_v_b_16')
// (6, 11, 'neigh_op_lft_2')
// (6, 11, 'sp4_v_b_5')
// (6, 12, 'neigh_op_bnl_2')

reg n213 = 0;
// (4, 10, 'neigh_op_tnr_4')
// (4, 11, 'neigh_op_rgt_4')
// (4, 12, 'neigh_op_bnr_4')
// (5, 10, 'neigh_op_top_4')
// (5, 11, 'lutff_4/out')
// (5, 12, 'neigh_op_bot_4')
// (6, 10, 'local_g2_4')
// (6, 10, 'lutff_2/in_0')
// (6, 10, 'neigh_op_tnl_4')
// (6, 11, 'neigh_op_lft_4')
// (6, 12, 'neigh_op_bnl_4')

reg n214 = 0;
// (4, 10, 'neigh_op_tnr_7')
// (4, 11, 'neigh_op_rgt_7')
// (4, 11, 'sp4_h_r_3')
// (4, 12, 'neigh_op_bnr_7')
// (5, 10, 'neigh_op_top_7')
// (5, 11, 'lutff_7/out')
// (5, 11, 'sp4_h_r_14')
// (5, 12, 'neigh_op_bot_7')
// (6, 10, 'neigh_op_tnl_7')
// (6, 11, 'neigh_op_lft_7')
// (6, 11, 'sp4_h_r_27')
// (6, 12, 'neigh_op_bnl_7')
// (7, 11, 'local_g2_6')
// (7, 11, 'lutff_6/in_0')
// (7, 11, 'sp4_h_r_38')
// (8, 11, 'sp4_h_l_38')

reg n215 = 0;
// (4, 10, 'sp4_h_r_7')
// (5, 10, 'local_g0_2')
// (5, 10, 'lutff_2/in_0')
// (5, 10, 'sp4_h_r_18')
// (6, 9, 'neigh_op_tnr_5')
// (6, 10, 'neigh_op_rgt_5')
// (6, 10, 'sp4_h_r_31')
// (6, 11, 'neigh_op_bnr_5')
// (7, 9, 'neigh_op_top_5')
// (7, 10, 'local_g0_5')
// (7, 10, 'lutff_5/out')
// (7, 10, 'lutff_6/in_1')
// (7, 10, 'sp4_h_r_42')
// (7, 11, 'neigh_op_bot_5')
// (8, 9, 'neigh_op_tnl_5')
// (8, 10, 'neigh_op_lft_5')
// (8, 10, 'sp4_h_l_42')
// (8, 11, 'neigh_op_bnl_5')

wire n216;
// (4, 11, 'neigh_op_tnr_0')
// (4, 12, 'neigh_op_rgt_0')
// (4, 13, 'neigh_op_bnr_0')
// (5, 0, 'span12_vert_23')
// (5, 1, 'sp12_v_b_23')
// (5, 2, 'sp12_v_b_20')
// (5, 3, 'sp12_v_b_19')
// (5, 4, 'sp12_v_b_16')
// (5, 5, 'sp12_v_b_15')
// (5, 6, 'sp12_v_b_12')
// (5, 7, 'sp12_v_b_11')
// (5, 8, 'sp12_v_b_8')
// (5, 9, 'local_g2_4')
// (5, 9, 'local_g2_7')
// (5, 9, 'lutff_0/in_2')
// (5, 9, 'lutff_4/in_2')
// (5, 9, 'lutff_6/in_3')
// (5, 9, 'sp12_v_b_7')
// (5, 9, 'sp4_r_v_b_36')
// (5, 10, 'sp12_v_b_4')
// (5, 10, 'sp4_r_v_b_25')
// (5, 11, 'local_g2_3')
// (5, 11, 'lutff_1/in_2')
// (5, 11, 'neigh_op_top_0')
// (5, 11, 'sp12_v_b_3')
// (5, 11, 'sp4_r_v_b_12')
// (5, 12, 'lutff_0/out')
// (5, 12, 'sp12_v_b_0')
// (5, 12, 'sp4_r_v_b_1')
// (5, 13, 'neigh_op_bot_0')
// (6, 8, 'sp4_v_t_36')
// (6, 9, 'sp4_v_b_36')
// (6, 10, 'sp4_v_b_25')
// (6, 11, 'neigh_op_tnl_0')
// (6, 11, 'sp4_v_b_12')
// (6, 12, 'neigh_op_lft_0')
// (6, 12, 'sp4_v_b_1')
// (6, 13, 'neigh_op_bnl_0')

reg n217 = 0;
// (4, 11, 'neigh_op_tnr_2')
// (4, 12, 'neigh_op_rgt_2')
// (4, 13, 'neigh_op_bnr_2')
// (5, 11, 'neigh_op_top_2')
// (5, 12, 'local_g1_2')
// (5, 12, 'lutff_2/out')
// (5, 12, 'lutff_3/in_0')
// (5, 13, 'neigh_op_bot_2')
// (6, 11, 'neigh_op_tnl_2')
// (6, 12, 'neigh_op_lft_2')
// (6, 13, 'neigh_op_bnl_2')

reg n218 = 0;
// (4, 11, 'neigh_op_tnr_3')
// (4, 12, 'neigh_op_rgt_3')
// (4, 13, 'neigh_op_bnr_3')
// (5, 11, 'neigh_op_top_3')
// (5, 12, 'lutff_3/out')
// (5, 13, 'local_g1_3')
// (5, 13, 'lutff_6/in_0')
// (5, 13, 'neigh_op_bot_3')
// (6, 11, 'neigh_op_tnl_3')
// (6, 12, 'neigh_op_lft_3')
// (6, 13, 'neigh_op_bnl_3')

reg n219 = 0;
// (4, 11, 'neigh_op_tnr_4')
// (4, 12, 'local_g3_4')
// (4, 12, 'lutff_7/in_0')
// (4, 12, 'neigh_op_rgt_4')
// (4, 13, 'neigh_op_bnr_4')
// (5, 11, 'neigh_op_top_4')
// (5, 12, 'lutff_4/out')
// (5, 13, 'neigh_op_bot_4')
// (6, 11, 'neigh_op_tnl_4')
// (6, 12, 'neigh_op_lft_4')
// (6, 13, 'neigh_op_bnl_4')

reg n220 = 0;
// (4, 11, 'neigh_op_tnr_5')
// (4, 12, 'neigh_op_rgt_5')
// (4, 13, 'neigh_op_bnr_5')
// (5, 5, 'sp12_v_t_22')
// (5, 6, 'sp12_v_b_22')
// (5, 7, 'sp12_v_b_21')
// (5, 8, 'sp12_v_b_18')
// (5, 9, 'sp12_v_b_17')
// (5, 10, 'sp12_v_b_14')
// (5, 11, 'local_g3_5')
// (5, 11, 'lutff_4/in_0')
// (5, 11, 'neigh_op_top_5')
// (5, 11, 'sp12_v_b_13')
// (5, 12, 'lutff_5/out')
// (5, 12, 'sp12_v_b_10')
// (5, 13, 'neigh_op_bot_5')
// (5, 13, 'sp12_v_b_9')
// (5, 14, 'sp12_v_b_6')
// (5, 15, 'sp12_v_b_5')
// (5, 16, 'sp12_v_b_2')
// (5, 17, 'span12_vert_1')
// (6, 11, 'neigh_op_tnl_5')
// (6, 12, 'neigh_op_lft_5')
// (6, 13, 'neigh_op_bnl_5')

reg n221 = 0;
// (4, 11, 'neigh_op_tnr_6')
// (4, 12, 'neigh_op_rgt_6')
// (4, 13, 'neigh_op_bnr_6')
// (5, 11, 'neigh_op_top_6')
// (5, 12, 'local_g0_6')
// (5, 12, 'lutff_4/in_0')
// (5, 12, 'lutff_6/out')
// (5, 13, 'neigh_op_bot_6')
// (6, 11, 'neigh_op_tnl_6')
// (6, 12, 'neigh_op_lft_6')
// (6, 13, 'neigh_op_bnl_6')

reg n222 = 0;
// (4, 11, 'neigh_op_tnr_7')
// (4, 12, 'neigh_op_rgt_7')
// (4, 13, 'neigh_op_bnr_7')
// (5, 11, 'neigh_op_top_7')
// (5, 12, 'local_g1_7')
// (5, 12, 'lutff_2/in_0')
// (5, 12, 'lutff_7/out')
// (5, 13, 'neigh_op_bot_7')
// (6, 11, 'neigh_op_tnl_7')
// (6, 12, 'neigh_op_lft_7')
// (6, 13, 'neigh_op_bnl_7')

wire \d_out[2] ;
// (4, 11, 'sp12_h_r_1')
// (5, 11, 'sp12_h_r_2')
// (6, 11, 'sp12_h_r_5')
// (7, 11, 'sp12_h_r_6')
// (8, 11, 'sp12_h_r_9')
// (9, 11, 'sp12_h_r_10')
// (10, 10, 'neigh_op_tnr_3')
// (10, 11, 'neigh_op_rgt_3')
// (10, 11, 'sp12_h_r_13')
// (10, 12, 'neigh_op_bnr_3')
// (11, 10, 'neigh_op_top_3')
// (11, 11, 'lutff_3/out')
// (11, 11, 'sp12_h_r_14')
// (11, 12, 'neigh_op_bot_3')
// (12, 10, 'neigh_op_tnl_3')
// (12, 11, 'neigh_op_lft_3')
// (12, 11, 'sp12_h_r_17')
// (12, 12, 'neigh_op_bnl_3')
// (13, 11, 'io_1/D_OUT_0')
// (13, 11, 'io_1/PAD')
// (13, 11, 'local_g0_1')
// (13, 11, 'span12_horz_17')

reg n224 = 0;
// (4, 11, 'sp4_h_r_1')
// (5, 11, 'local_g1_4')
// (5, 11, 'lutff_6/in_1')
// (5, 11, 'sp4_h_r_12')
// (6, 10, 'neigh_op_tnr_2')
// (6, 11, 'neigh_op_rgt_2')
// (6, 11, 'sp4_h_r_25')
// (6, 12, 'neigh_op_bnr_2')
// (7, 10, 'neigh_op_top_2')
// (7, 11, 'local_g2_2')
// (7, 11, 'lutff_0/in_0')
// (7, 11, 'lutff_2/out')
// (7, 11, 'sp4_h_r_36')
// (7, 12, 'neigh_op_bot_2')
// (8, 10, 'neigh_op_tnl_2')
// (8, 11, 'neigh_op_lft_2')
// (8, 11, 'sp4_h_l_36')
// (8, 12, 'neigh_op_bnl_2')

reg n225 = 0;
// (4, 11, 'sp4_r_v_b_39')
// (4, 12, 'sp4_r_v_b_26')
// (4, 13, 'neigh_op_tnr_1')
// (4, 13, 'sp4_r_v_b_15')
// (4, 14, 'neigh_op_rgt_1')
// (4, 14, 'sp4_r_v_b_2')
// (4, 15, 'neigh_op_bnr_1')
// (5, 10, 'sp4_v_t_39')
// (5, 11, 'sp4_v_b_39')
// (5, 12, 'local_g3_2')
// (5, 12, 'lutff_7/in_0')
// (5, 12, 'sp4_v_b_26')
// (5, 13, 'local_g0_1')
// (5, 13, 'local_g1_1')
// (5, 13, 'lutff_0/in_0')
// (5, 13, 'lutff_7/in_0')
// (5, 13, 'neigh_op_top_1')
// (5, 13, 'sp4_v_b_15')
// (5, 14, 'local_g1_1')
// (5, 14, 'lutff_1/out')
// (5, 14, 'lutff_4/in_0')
// (5, 14, 'sp4_v_b_2')
// (5, 15, 'neigh_op_bot_1')
// (6, 13, 'neigh_op_tnl_1')
// (6, 14, 'neigh_op_lft_1')
// (6, 15, 'neigh_op_bnl_1')

wire n226;
// (4, 12, 'neigh_op_tnr_0')
// (4, 13, 'neigh_op_rgt_0')
// (4, 14, 'neigh_op_bnr_0')
// (5, 12, 'local_g1_0')
// (5, 12, 'lutff_0/in_3')
// (5, 12, 'neigh_op_top_0')
// (5, 13, 'lutff_0/out')
// (5, 14, 'neigh_op_bot_0')
// (6, 12, 'neigh_op_tnl_0')
// (6, 13, 'neigh_op_lft_0')
// (6, 14, 'neigh_op_bnl_0')

wire n227;
// (4, 12, 'neigh_op_tnr_1')
// (4, 13, 'neigh_op_rgt_1')
// (4, 14, 'neigh_op_bnr_1')
// (5, 12, 'neigh_op_top_1')
// (5, 13, 'local_g2_1')
// (5, 13, 'lutff_0/in_3')
// (5, 13, 'lutff_1/out')
// (5, 14, 'neigh_op_bot_1')
// (6, 12, 'neigh_op_tnl_1')
// (6, 13, 'neigh_op_lft_1')
// (6, 14, 'neigh_op_bnl_1')

reg n228 = 0;
// (4, 12, 'neigh_op_tnr_2')
// (4, 13, 'neigh_op_rgt_2')
// (4, 14, 'neigh_op_bnr_2')
// (5, 12, 'neigh_op_top_2')
// (5, 13, 'local_g1_2')
// (5, 13, 'lutff_1/in_0')
// (5, 13, 'lutff_2/out')
// (5, 14, 'local_g1_2')
// (5, 14, 'lutff_4/in_1')
// (5, 14, 'neigh_op_bot_2')
// (6, 12, 'neigh_op_tnl_2')
// (6, 13, 'neigh_op_lft_2')
// (6, 14, 'neigh_op_bnl_2')

reg n229 = 0;
// (4, 12, 'neigh_op_tnr_5')
// (4, 13, 'neigh_op_rgt_5')
// (4, 14, 'neigh_op_bnr_5')
// (5, 12, 'neigh_op_top_5')
// (5, 13, 'local_g0_5')
// (5, 13, 'lutff_3/in_0')
// (5, 13, 'lutff_5/out')
// (5, 14, 'neigh_op_bot_5')
// (6, 12, 'neigh_op_tnl_5')
// (6, 13, 'neigh_op_lft_5')
// (6, 14, 'neigh_op_bnl_5')

reg n230 = 0;
// (4, 12, 'neigh_op_tnr_6')
// (4, 13, 'neigh_op_rgt_6')
// (4, 14, 'neigh_op_bnr_6')
// (5, 12, 'neigh_op_top_6')
// (5, 13, 'local_g2_6')
// (5, 13, 'lutff_1/in_1')
// (5, 13, 'lutff_6/out')
// (5, 13, 'lutff_7/in_1')
// (5, 14, 'neigh_op_bot_6')
// (6, 12, 'neigh_op_tnl_6')
// (6, 13, 'neigh_op_lft_6')
// (6, 14, 'neigh_op_bnl_6')

reg n231 = 0;
// (4, 12, 'neigh_op_tnr_7')
// (4, 13, 'neigh_op_rgt_7')
// (4, 14, 'neigh_op_bnr_7')
// (5, 12, 'neigh_op_top_7')
// (5, 13, 'local_g0_7')
// (5, 13, 'lutff_5/in_0')
// (5, 13, 'lutff_7/out')
// (5, 14, 'neigh_op_bot_7')
// (6, 12, 'neigh_op_tnl_7')
// (6, 13, 'neigh_op_lft_7')
// (6, 14, 'neigh_op_bnl_7')

reg n232 = 0;
// (4, 13, 'neigh_op_tnr_3')
// (4, 14, 'neigh_op_rgt_3')
// (4, 15, 'neigh_op_bnr_3')
// (5, 13, 'neigh_op_top_3')
// (5, 14, 'local_g0_3')
// (5, 14, 'lutff_3/out')
// (5, 14, 'lutff_7/in_0')
// (5, 15, 'neigh_op_bot_3')
// (6, 13, 'neigh_op_tnl_3')
// (6, 14, 'neigh_op_lft_3')
// (6, 15, 'neigh_op_bnl_3')

reg n233 = 0;
// (4, 13, 'neigh_op_tnr_4')
// (4, 14, 'neigh_op_rgt_4')
// (4, 15, 'neigh_op_bnr_4')
// (5, 13, 'neigh_op_top_4')
// (5, 14, 'local_g1_4')
// (5, 14, 'lutff_3/in_0')
// (5, 14, 'lutff_4/out')
// (5, 15, 'neigh_op_bot_4')
// (6, 13, 'neigh_op_tnl_4')
// (6, 14, 'neigh_op_lft_4')
// (6, 15, 'neigh_op_bnl_4')

reg n234 = 0;
// (4, 13, 'neigh_op_tnr_5')
// (4, 14, 'neigh_op_rgt_5')
// (4, 15, 'neigh_op_bnr_5')
// (5, 13, 'neigh_op_top_5')
// (5, 14, 'lutff_5/out')
// (5, 15, 'neigh_op_bot_5')
// (6, 13, 'neigh_op_tnl_5')
// (6, 14, 'local_g1_5')
// (6, 14, 'lutff_2/in_0')
// (6, 14, 'neigh_op_lft_5')
// (6, 15, 'neigh_op_bnl_5')

reg n235 = 0;
// (4, 13, 'neigh_op_tnr_7')
// (4, 14, 'neigh_op_rgt_7')
// (4, 15, 'neigh_op_bnr_7')
// (5, 13, 'neigh_op_top_7')
// (5, 14, 'local_g0_7')
// (5, 14, 'lutff_1/in_0')
// (5, 14, 'lutff_7/out')
// (5, 15, 'neigh_op_bot_7')
// (6, 13, 'neigh_op_tnl_7')
// (6, 14, 'neigh_op_lft_7')
// (6, 15, 'neigh_op_bnl_7')

wire n236;
// (5, 1, 'neigh_op_tnr_1')
// (5, 2, 'neigh_op_rgt_1')
// (5, 3, 'neigh_op_bnr_1')
// (6, 1, 'neigh_op_top_1')
// (6, 1, 'sp4_r_v_b_14')
// (6, 2, 'lutff_1/out')
// (6, 2, 'sp4_r_v_b_3')
// (6, 3, 'neigh_op_bot_1')
// (6, 3, 'sp4_r_v_b_43')
// (6, 4, 'sp4_r_v_b_30')
// (6, 5, 'sp4_r_v_b_19')
// (6, 6, 'sp4_r_v_b_6')
// (7, 0, 'span4_vert_14')
// (7, 1, 'neigh_op_tnl_1')
// (7, 1, 'sp4_v_b_14')
// (7, 2, 'neigh_op_lft_1')
// (7, 2, 'sp4_v_b_3')
// (7, 2, 'sp4_v_t_43')
// (7, 3, 'local_g2_3')
// (7, 3, 'lutff_2/in_3')
// (7, 3, 'lutff_6/in_3')
// (7, 3, 'neigh_op_bnl_1')
// (7, 3, 'sp4_v_b_43')
// (7, 4, 'sp4_v_b_30')
// (7, 5, 'sp4_v_b_19')
// (7, 6, 'sp4_v_b_6')

wire n237;
// (5, 1, 'neigh_op_tnr_2')
// (5, 2, 'neigh_op_rgt_2')
// (5, 3, 'neigh_op_bnr_2')
// (6, 1, 'neigh_op_top_2')
// (6, 2, 'lutff_2/out')
// (6, 2, 'sp4_r_v_b_37')
// (6, 3, 'local_g1_0')
// (6, 3, 'lutff_4/in_3')
// (6, 3, 'neigh_op_bot_2')
// (6, 3, 'sp4_r_v_b_24')
// (6, 4, 'sp4_r_v_b_13')
// (6, 5, 'sp4_r_v_b_0')
// (7, 1, 'neigh_op_tnl_2')
// (7, 1, 'sp4_v_t_37')
// (7, 2, 'neigh_op_lft_2')
// (7, 2, 'sp4_v_b_37')
// (7, 3, 'local_g2_2')
// (7, 3, 'lutff_1/in_3')
// (7, 3, 'neigh_op_bnl_2')
// (7, 3, 'sp4_v_b_24')
// (7, 4, 'sp4_v_b_13')
// (7, 5, 'sp4_v_b_0')

wire n238;
// (5, 1, 'neigh_op_tnr_3')
// (5, 2, 'neigh_op_rgt_3')
// (5, 3, 'neigh_op_bnr_3')
// (6, 1, 'neigh_op_top_3')
// (6, 2, 'local_g0_3')
// (6, 2, 'local_g1_3')
// (6, 2, 'lutff_1/in_0')
// (6, 2, 'lutff_2/in_0')
// (6, 2, 'lutff_3/out')
// (6, 3, 'local_g0_3')
// (6, 3, 'lutff_5/in_2')
// (6, 3, 'neigh_op_bot_3')
// (7, 1, 'neigh_op_tnl_3')
// (7, 2, 'neigh_op_lft_3')
// (7, 3, 'neigh_op_bnl_3')

wire n239;
// (5, 1, 'neigh_op_tnr_5')
// (5, 2, 'neigh_op_rgt_5')
// (5, 3, 'neigh_op_bnr_5')
// (6, 1, 'neigh_op_top_5')
// (6, 2, 'lutff_5/out')
// (6, 3, 'local_g0_5')
// (6, 3, 'local_g1_5')
// (6, 3, 'lutff_0/in_0')
// (6, 3, 'lutff_1/in_1')
// (6, 3, 'lutff_2/in_3')
// (6, 3, 'lutff_3/in_2')
// (6, 3, 'lutff_5/in_1')
// (6, 3, 'lutff_6/in_2')
// (6, 3, 'lutff_7/in_0')
// (6, 3, 'neigh_op_bot_5')
// (7, 1, 'neigh_op_tnl_5')
// (7, 2, 'neigh_op_lft_5')
// (7, 3, 'neigh_op_bnl_5')

wire n240;
// (5, 1, 'neigh_op_tnr_6')
// (5, 2, 'neigh_op_rgt_6')
// (5, 3, 'neigh_op_bnr_6')
// (6, 1, 'neigh_op_top_6')
// (6, 2, 'local_g0_6')
// (6, 2, 'local_g1_6')
// (6, 2, 'lutff_3/in_1')
// (6, 2, 'lutff_5/in_2')
// (6, 2, 'lutff_6/out')
// (6, 3, 'neigh_op_bot_6')
// (7, 1, 'neigh_op_tnl_6')
// (7, 2, 'neigh_op_lft_6')
// (7, 3, 'neigh_op_bnl_6')

wire n241;
// (5, 1, 'neigh_op_tnr_7')
// (5, 2, 'neigh_op_rgt_7')
// (5, 3, 'neigh_op_bnr_7')
// (6, 1, 'neigh_op_top_7')
// (6, 2, 'local_g0_7')
// (6, 2, 'lutff_2/in_3')
// (6, 2, 'lutff_7/out')
// (6, 3, 'neigh_op_bot_7')
// (7, 1, 'neigh_op_tnl_7')
// (7, 2, 'neigh_op_lft_7')
// (7, 3, 'neigh_op_bnl_7')

wire n242;
// (5, 1, 'sp4_r_v_b_42')
// (5, 2, 'sp4_h_r_9')
// (5, 2, 'sp4_r_v_b_31')
// (5, 3, 'sp4_r_v_b_18')
// (5, 4, 'sp4_r_v_b_7')
// (6, 0, 'span4_vert_42')
// (6, 1, 'sp4_v_b_42')
// (6, 2, 'local_g0_4')
// (6, 2, 'local_g1_4')
// (6, 2, 'lutff_6/in_3')
// (6, 2, 'lutff_7/in_3')
// (6, 2, 'sp4_h_r_20')
// (6, 2, 'sp4_v_b_31')
// (6, 3, 'local_g0_2')
// (6, 3, 'lutff_4/in_2')
// (6, 3, 'sp4_v_b_18')
// (6, 4, 'sp4_h_r_2')
// (6, 4, 'sp4_v_b_7')
// (7, 1, 'sp4_r_v_b_47')
// (7, 2, 'local_g2_1')
// (7, 2, 'local_g2_2')
// (7, 2, 'lutff_3/in_2')
// (7, 2, 'lutff_7/in_3')
// (7, 2, 'sp4_h_r_33')
// (7, 2, 'sp4_r_v_b_34')
// (7, 3, 'neigh_op_tnr_5')
// (7, 3, 'sp4_r_v_b_23')
// (7, 4, 'neigh_op_rgt_5')
// (7, 4, 'sp4_h_r_15')
// (7, 4, 'sp4_r_v_b_10')
// (7, 5, 'neigh_op_bnr_5')
// (8, 0, 'span4_vert_47')
// (8, 1, 'sp4_v_b_47')
// (8, 2, 'sp4_h_r_44')
// (8, 2, 'sp4_v_b_34')
// (8, 3, 'neigh_op_top_5')
// (8, 3, 'sp4_r_v_b_38')
// (8, 3, 'sp4_v_b_23')
// (8, 4, 'lutff_5/out')
// (8, 4, 'sp4_h_r_26')
// (8, 4, 'sp4_r_v_b_27')
// (8, 4, 'sp4_v_b_10')
// (8, 5, 'neigh_op_bot_5')
// (8, 5, 'sp4_r_v_b_14')
// (8, 6, 'sp4_r_v_b_3')
// (9, 2, 'sp4_h_l_44')
// (9, 2, 'sp4_v_t_38')
// (9, 3, 'neigh_op_tnl_5')
// (9, 3, 'sp4_v_b_38')
// (9, 4, 'neigh_op_lft_5')
// (9, 4, 'sp4_h_r_39')
// (9, 4, 'sp4_v_b_27')
// (9, 5, 'neigh_op_bnl_5')
// (9, 5, 'sp4_v_b_14')
// (9, 6, 'sp4_v_b_3')
// (10, 4, 'sp4_h_l_39')

wire n243;
// (5, 2, 'neigh_op_tnr_2')
// (5, 3, 'neigh_op_rgt_2')
// (5, 4, 'neigh_op_bnr_2')
// (6, 2, 'neigh_op_top_2')
// (6, 3, 'local_g1_2')
// (6, 3, 'lutff_2/out')
// (6, 3, 'lutff_4/in_1')
// (6, 3, 'sp4_h_r_4')
// (6, 4, 'neigh_op_bot_2')
// (7, 2, 'neigh_op_tnl_2')
// (7, 3, 'local_g1_1')
// (7, 3, 'lutff_2/in_0')
// (7, 3, 'neigh_op_lft_2')
// (7, 3, 'sp4_h_r_17')
// (7, 4, 'neigh_op_bnl_2')
// (8, 3, 'sp4_h_r_28')
// (9, 3, 'sp4_h_r_41')
// (10, 3, 'sp4_h_l_41')

wire n244;
// (5, 2, 'neigh_op_tnr_3')
// (5, 3, 'neigh_op_rgt_3')
// (5, 3, 'sp4_h_r_11')
// (5, 4, 'neigh_op_bnr_3')
// (6, 2, 'neigh_op_top_3')
// (6, 3, 'lutff_3/out')
// (6, 3, 'sp4_h_r_22')
// (6, 4, 'neigh_op_bot_3')
// (7, 2, 'neigh_op_tnl_3')
// (7, 3, 'neigh_op_lft_3')
// (7, 3, 'sp4_h_r_35')
// (7, 4, 'local_g3_3')
// (7, 4, 'lutff_0/in_0')
// (7, 4, 'neigh_op_bnl_3')
// (8, 3, 'local_g2_6')
// (8, 3, 'lutff_0/in_0')
// (8, 3, 'sp4_h_r_46')
// (9, 3, 'sp4_h_l_46')

wire n245;
// (5, 2, 'neigh_op_tnr_4')
// (5, 3, 'neigh_op_rgt_4')
// (5, 3, 'sp4_r_v_b_40')
// (5, 4, 'neigh_op_bnr_4')
// (5, 4, 'sp4_r_v_b_29')
// (5, 5, 'sp4_r_v_b_16')
// (5, 6, 'sp4_r_v_b_5')
// (6, 1, 'sp4_r_v_b_33')
// (6, 2, 'neigh_op_top_4')
// (6, 2, 'sp4_r_v_b_20')
// (6, 2, 'sp4_v_t_40')
// (6, 3, 'lutff_4/out')
// (6, 3, 'sp4_r_v_b_9')
// (6, 3, 'sp4_v_b_40')
// (6, 4, 'local_g0_4')
// (6, 4, 'local_g2_5')
// (6, 4, 'lutff_1/in_2')
// (6, 4, 'lutff_7/in_1')
// (6, 4, 'neigh_op_bot_4')
// (6, 4, 'sp4_v_b_29')
// (6, 5, 'sp4_v_b_16')
// (6, 6, 'sp4_v_b_5')
// (7, 0, 'span4_vert_33')
// (7, 1, 'sp4_v_b_33')
// (7, 2, 'neigh_op_tnl_4')
// (7, 2, 'sp4_v_b_20')
// (7, 3, 'local_g0_1')
// (7, 3, 'lutff_5/in_0')
// (7, 3, 'neigh_op_lft_4')
// (7, 3, 'sp4_v_b_9')
// (7, 4, 'neigh_op_bnl_4')

wire n246;
// (5, 2, 'neigh_op_tnr_6')
// (5, 3, 'neigh_op_rgt_6')
// (5, 4, 'neigh_op_bnr_6')
// (6, 2, 'neigh_op_top_6')
// (6, 3, 'lutff_6/out')
// (6, 4, 'neigh_op_bot_6')
// (7, 2, 'neigh_op_tnl_6')
// (7, 3, 'local_g0_6')
// (7, 3, 'local_g1_6')
// (7, 3, 'lutff_0/in_1')
// (7, 3, 'lutff_3/in_1')
// (7, 3, 'lutff_4/in_1')
// (7, 3, 'lutff_7/in_2')
// (7, 3, 'neigh_op_lft_6')
// (7, 4, 'neigh_op_bnl_6')

wire n247;
// (5, 2, 'neigh_op_tnr_7')
// (5, 3, 'neigh_op_rgt_7')
// (5, 4, 'neigh_op_bnr_7')
// (6, 2, 'neigh_op_top_7')
// (6, 3, 'lutff_7/out')
// (6, 4, 'neigh_op_bot_7')
// (7, 2, 'neigh_op_tnl_7')
// (7, 3, 'local_g0_7')
// (7, 3, 'local_g1_7')
// (7, 3, 'lutff_0/in_0')
// (7, 3, 'lutff_3/in_0')
// (7, 3, 'lutff_4/in_0')
// (7, 3, 'lutff_7/in_0')
// (7, 3, 'neigh_op_lft_7')
// (7, 4, 'neigh_op_bnl_7')

wire n248;
// (5, 2, 'sp4_h_r_4')
// (6, 2, 'local_g0_1')
// (6, 2, 'local_g1_1')
// (6, 2, 'lutff_6/in_2')
// (6, 2, 'lutff_7/in_2')
// (6, 2, 'sp4_h_r_17')
// (7, 1, 'neigh_op_tnr_5')
// (7, 2, 'local_g3_5')
// (7, 2, 'lutff_3/in_1')
// (7, 2, 'neigh_op_rgt_5')
// (7, 2, 'sp4_h_r_28')
// (7, 3, 'local_g0_5')
// (7, 3, 'lutff_1/in_0')
// (7, 3, 'neigh_op_bnr_5')
// (8, 1, 'neigh_op_top_5')
// (8, 1, 'sp4_r_v_b_22')
// (8, 2, 'lutff_5/out')
// (8, 2, 'sp4_h_r_41')
// (8, 2, 'sp4_r_v_b_11')
// (8, 3, 'neigh_op_bot_5')
// (9, 0, 'span4_vert_22')
// (9, 1, 'neigh_op_tnl_5')
// (9, 1, 'sp4_v_b_22')
// (9, 2, 'neigh_op_lft_5')
// (9, 2, 'sp4_h_l_41')
// (9, 2, 'sp4_v_b_11')
// (9, 3, 'neigh_op_bnl_5')

wire n249;
// (5, 3, 'neigh_op_tnr_0')
// (5, 4, 'neigh_op_rgt_0')
// (5, 5, 'neigh_op_bnr_0')
// (6, 3, 'neigh_op_top_0')
// (6, 4, 'local_g0_0')
// (6, 4, 'lutff_0/out')
// (6, 4, 'lutff_1/in_1')
// (6, 5, 'neigh_op_bot_0')
// (7, 3, 'neigh_op_tnl_0')
// (7, 4, 'neigh_op_lft_0')
// (7, 5, 'neigh_op_bnl_0')

wire n250;
// (5, 3, 'neigh_op_tnr_1')
// (5, 4, 'neigh_op_rgt_1')
// (5, 5, 'neigh_op_bnr_1')
// (6, 3, 'neigh_op_top_1')
// (6, 4, 'lutff_1/out')
// (6, 5, 'neigh_op_bot_1')
// (7, 3, 'neigh_op_tnl_1')
// (7, 4, 'local_g0_1')
// (7, 4, 'lutff_4/in_1')
// (7, 4, 'neigh_op_lft_1')
// (7, 5, 'neigh_op_bnl_1')

wire n251;
// (5, 3, 'neigh_op_tnr_2')
// (5, 4, 'neigh_op_rgt_2')
// (5, 5, 'neigh_op_bnr_2')
// (6, 3, 'neigh_op_top_2')
// (6, 4, 'local_g2_2')
// (6, 4, 'lutff_2/out')
// (6, 4, 'lutff_7/in_3')
// (6, 5, 'neigh_op_bot_2')
// (7, 3, 'neigh_op_tnl_2')
// (7, 4, 'neigh_op_lft_2')
// (7, 5, 'neigh_op_bnl_2')

wire n252;
// (5, 3, 'neigh_op_tnr_4')
// (5, 4, 'neigh_op_rgt_4')
// (5, 5, 'neigh_op_bnr_4')
// (6, 3, 'neigh_op_top_4')
// (6, 4, 'local_g1_4')
// (6, 4, 'lutff_1/in_0')
// (6, 4, 'lutff_4/out')
// (6, 5, 'local_g1_4')
// (6, 5, 'lutff_3/in_2')
// (6, 5, 'neigh_op_bot_4')
// (7, 3, 'neigh_op_tnl_4')
// (7, 4, 'neigh_op_lft_4')
// (7, 5, 'neigh_op_bnl_4')

wire n253;
// (5, 3, 'neigh_op_tnr_7')
// (5, 4, 'neigh_op_rgt_7')
// (5, 5, 'neigh_op_bnr_7')
// (6, 2, 'sp4_r_v_b_39')
// (6, 3, 'neigh_op_top_7')
// (6, 3, 'sp4_r_v_b_26')
// (6, 4, 'lutff_7/out')
// (6, 4, 'sp4_r_v_b_15')
// (6, 5, 'neigh_op_bot_7')
// (6, 5, 'sp4_r_v_b_2')
// (7, 1, 'sp4_v_t_39')
// (7, 2, 'sp4_v_b_39')
// (7, 3, 'neigh_op_tnl_7')
// (7, 3, 'sp4_v_b_26')
// (7, 4, 'neigh_op_lft_7')
// (7, 4, 'sp4_v_b_15')
// (7, 5, 'neigh_op_bnl_7')
// (7, 5, 'sp4_h_r_8')
// (7, 5, 'sp4_v_b_2')
// (8, 5, 'local_g1_5')
// (8, 5, 'lutff_2/in_2')
// (8, 5, 'sp4_h_r_21')
// (9, 5, 'sp4_h_r_32')
// (10, 5, 'sp4_h_r_45')
// (11, 5, 'sp4_h_l_45')

wire n254;
// (5, 3, 'sp4_h_r_3')
// (6, 2, 'sp4_h_r_5')
// (6, 3, 'sp4_h_r_14')
// (7, 2, 'local_g0_0')
// (7, 2, 'lutff_0/in_2')
// (7, 2, 'sp4_h_r_16')
// (7, 3, 'local_g3_3')
// (7, 3, 'lutff_6/in_2')
// (7, 3, 'sp4_h_r_27')
// (8, 2, 'local_g2_5')
// (8, 2, 'lutff_3/in_2')
// (8, 2, 'sp4_h_r_29')
// (8, 3, 'neigh_op_tnr_6')
// (8, 3, 'sp4_h_r_38')
// (8, 4, 'neigh_op_rgt_6')
// (8, 4, 'sp4_r_v_b_44')
// (8, 5, 'neigh_op_bnr_6')
// (8, 5, 'sp4_r_v_b_33')
// (8, 6, 'sp4_r_v_b_20')
// (8, 7, 'sp4_r_v_b_9')
// (9, 2, 'sp4_h_r_40')
// (9, 3, 'neigh_op_top_6')
// (9, 3, 'sp4_h_l_38')
// (9, 3, 'sp4_h_r_2')
// (9, 3, 'sp4_r_v_b_40')
// (9, 3, 'sp4_v_t_44')
// (9, 4, 'lutff_6/out')
// (9, 4, 'sp4_r_v_b_29')
// (9, 4, 'sp4_v_b_44')
// (9, 5, 'neigh_op_bot_6')
// (9, 5, 'sp4_r_v_b_16')
// (9, 5, 'sp4_v_b_33')
// (9, 6, 'sp4_r_v_b_5')
// (9, 6, 'sp4_v_b_20')
// (9, 7, 'sp4_v_b_9')
// (10, 2, 'sp4_h_l_40')
// (10, 2, 'sp4_v_t_40')
// (10, 3, 'neigh_op_tnl_6')
// (10, 3, 'sp4_h_r_15')
// (10, 3, 'sp4_v_b_40')
// (10, 4, 'neigh_op_lft_6')
// (10, 4, 'sp4_v_b_29')
// (10, 5, 'neigh_op_bnl_6')
// (10, 5, 'sp4_v_b_16')
// (10, 6, 'sp4_v_b_5')
// (11, 3, 'local_g2_2')
// (11, 3, 'lutff_5/in_3')
// (11, 3, 'sp4_h_r_26')
// (12, 3, 'sp4_h_r_39')
// (13, 3, 'span4_horz_39')

wire n255;
// (5, 4, 'neigh_op_tnr_1')
// (5, 5, 'local_g2_1')
// (5, 5, 'local_g3_1')
// (5, 5, 'lutff_2/in_2')
// (5, 5, 'lutff_7/in_2')
// (5, 5, 'neigh_op_rgt_1')
// (5, 6, 'neigh_op_bnr_1')
// (6, 2, 'sp12_v_t_22')
// (6, 3, 'sp12_v_b_22')
// (6, 4, 'neigh_op_top_1')
// (6, 4, 'sp12_v_b_21')
// (6, 4, 'sp4_r_v_b_46')
// (6, 5, 'lutff_1/out')
// (6, 5, 'sp12_v_b_18')
// (6, 5, 'sp4_r_v_b_35')
// (6, 6, 'neigh_op_bot_1')
// (6, 6, 'sp12_v_b_17')
// (6, 6, 'sp4_r_v_b_22')
// (6, 7, 'local_g2_3')
// (6, 7, 'lutff_7/in_0')
// (6, 7, 'sp12_v_b_14')
// (6, 7, 'sp4_r_v_b_11')
// (6, 8, 'local_g3_5')
// (6, 8, 'lutff_6/in_2')
// (6, 8, 'sp12_v_b_13')
// (6, 9, 'sp12_v_b_10')
// (6, 10, 'sp12_v_b_9')
// (6, 11, 'sp12_v_b_6')
// (6, 12, 'sp12_v_b_5')
// (6, 13, 'sp12_v_b_2')
// (6, 14, 'sp12_v_b_1')
// (7, 3, 'sp4_v_t_46')
// (7, 4, 'neigh_op_tnl_1')
// (7, 4, 'sp4_v_b_46')
// (7, 5, 'neigh_op_lft_1')
// (7, 5, 'sp4_v_b_35')
// (7, 6, 'neigh_op_bnl_1')
// (7, 6, 'sp4_v_b_22')
// (7, 7, 'sp4_v_b_11')

wire n256;
// (5, 4, 'neigh_op_tnr_2')
// (5, 5, 'neigh_op_rgt_2')
// (5, 6, 'neigh_op_bnr_2')
// (6, 4, 'neigh_op_top_2')
// (6, 5, 'local_g1_2')
// (6, 5, 'lutff_1/in_2')
// (6, 5, 'lutff_2/out')
// (6, 6, 'neigh_op_bot_2')
// (7, 4, 'neigh_op_tnl_2')
// (7, 5, 'neigh_op_lft_2')
// (7, 6, 'neigh_op_bnl_2')

wire n257;
// (5, 4, 'neigh_op_tnr_3')
// (5, 5, 'neigh_op_rgt_3')
// (5, 6, 'neigh_op_bnr_3')
// (6, 4, 'neigh_op_top_3')
// (6, 5, 'lutff_3/out')
// (6, 6, 'neigh_op_bot_3')
// (7, 4, 'neigh_op_tnl_3')
// (7, 5, 'local_g0_3')
// (7, 5, 'lutff_5/in_2')
// (7, 5, 'neigh_op_lft_3')
// (7, 6, 'neigh_op_bnl_3')

wire n258;
// (5, 4, 'neigh_op_tnr_4')
// (5, 5, 'neigh_op_rgt_4')
// (5, 6, 'neigh_op_bnr_4')
// (6, 4, 'neigh_op_top_4')
// (6, 5, 'lutff_4/out')
// (6, 6, 'neigh_op_bot_4')
// (7, 4, 'neigh_op_tnl_4')
// (7, 5, 'local_g0_4')
// (7, 5, 'lutff_2/in_2')
// (7, 5, 'neigh_op_lft_4')
// (7, 6, 'neigh_op_bnl_4')

wire n259;
// (5, 4, 'neigh_op_tnr_5')
// (5, 5, 'neigh_op_rgt_5')
// (5, 6, 'neigh_op_bnr_5')
// (6, 4, 'neigh_op_top_5')
// (6, 5, 'lutff_5/out')
// (6, 6, 'neigh_op_bot_5')
// (7, 4, 'neigh_op_tnl_5')
// (7, 5, 'local_g1_5')
// (7, 5, 'lutff_0/in_2')
// (7, 5, 'neigh_op_lft_5')
// (7, 6, 'neigh_op_bnl_5')

wire n260;
// (5, 4, 'neigh_op_tnr_6')
// (5, 5, 'neigh_op_rgt_6')
// (5, 6, 'neigh_op_bnr_6')
// (6, 4, 'neigh_op_top_6')
// (6, 5, 'local_g0_6')
// (6, 5, 'lutff_2/in_2')
// (6, 5, 'lutff_4/in_0')
// (6, 5, 'lutff_6/out')
// (6, 6, 'neigh_op_bot_6')
// (7, 4, 'neigh_op_tnl_6')
// (7, 5, 'neigh_op_lft_6')
// (7, 6, 'neigh_op_bnl_6')

reg n261 = 0;
// (5, 4, 'neigh_op_tnr_7')
// (5, 5, 'local_g2_7')
// (5, 5, 'lutff_3/in_0')
// (5, 5, 'neigh_op_rgt_7')
// (5, 6, 'neigh_op_bnr_7')
// (6, 4, 'neigh_op_top_7')
// (6, 5, 'lutff_7/out')
// (6, 6, 'neigh_op_bot_7')
// (7, 4, 'neigh_op_tnl_7')
// (7, 5, 'neigh_op_lft_7')
// (7, 6, 'neigh_op_bnl_7')

wire n262;
// (5, 4, 'sp12_h_r_1')
// (6, 4, 'sp12_h_r_2')
// (7, 3, 'neigh_op_tnr_7')
// (7, 3, 'sp4_r_v_b_43')
// (7, 4, 'neigh_op_rgt_7')
// (7, 4, 'sp12_h_r_5')
// (7, 4, 'sp4_r_v_b_30')
// (7, 5, 'neigh_op_bnr_7')
// (7, 5, 'sp4_r_v_b_19')
// (7, 6, 'sp4_r_v_b_6')
// (7, 7, 'sp4_r_v_b_44')
// (7, 8, 'sp4_r_v_b_33')
// (7, 9, 'sp4_r_v_b_20')
// (7, 10, 'sp4_r_v_b_9')
// (8, 0, 'span12_vert_21')
// (8, 1, 'sp12_v_b_21')
// (8, 2, 'sp12_v_b_18')
// (8, 2, 'sp4_v_t_43')
// (8, 3, 'neigh_op_top_7')
// (8, 3, 'sp12_v_b_17')
// (8, 3, 'sp4_v_b_43')
// (8, 4, 'lutff_7/out')
// (8, 4, 'sp12_h_r_6')
// (8, 4, 'sp12_v_b_14')
// (8, 4, 'sp4_v_b_30')
// (8, 5, 'neigh_op_bot_7')
// (8, 5, 'sp12_v_b_13')
// (8, 5, 'sp4_v_b_19')
// (8, 6, 'sp12_v_b_10')
// (8, 6, 'sp4_v_b_6')
// (8, 6, 'sp4_v_t_44')
// (8, 7, 'sp12_v_b_9')
// (8, 7, 'sp4_v_b_44')
// (8, 8, 'sp12_v_b_6')
// (8, 8, 'sp4_v_b_33')
// (8, 9, 'local_g0_4')
// (8, 9, 'lutff_6/in_2')
// (8, 9, 'sp12_v_b_5')
// (8, 9, 'sp4_v_b_20')
// (8, 10, 'sp12_v_b_2')
// (8, 10, 'sp4_v_b_9')
// (8, 11, 'sp12_h_r_1')
// (8, 11, 'sp12_v_b_1')
// (9, 3, 'neigh_op_tnl_7')
// (9, 4, 'neigh_op_lft_7')
// (9, 4, 'sp12_h_r_9')
// (9, 5, 'neigh_op_bnl_7')
// (9, 11, 'sp12_h_r_2')
// (10, 4, 'sp12_h_r_10')
// (10, 11, 'sp12_h_r_5')
// (11, 4, 'local_g0_5')
// (11, 4, 'lutff_7/in_0')
// (11, 4, 'sp12_h_r_13')
// (11, 11, 'local_g0_6')
// (11, 11, 'local_g1_6')
// (11, 11, 'lutff_1/in_2')
// (11, 11, 'lutff_4/in_2')
// (11, 11, 'sp12_h_r_6')
// (12, 4, 'sp12_h_r_14')
// (12, 11, 'sp12_h_r_9')
// (13, 4, 'span12_horz_14')
// (13, 11, 'span12_horz_9')

wire n263;
// (5, 4, 'sp4_r_v_b_39')
// (5, 4, 'sp4_r_v_b_43')
// (5, 5, 'sp4_r_v_b_26')
// (5, 5, 'sp4_r_v_b_30')
// (5, 6, 'local_g2_7')
// (5, 6, 'local_g3_1')
// (5, 6, 'lutff_4/in_1')
// (5, 6, 'lutff_5/in_3')
// (5, 6, 'sp4_r_v_b_15')
// (5, 6, 'sp4_r_v_b_19')
// (5, 6, 'sp4_r_v_b_41')
// (5, 7, 'local_g0_4')
// (5, 7, 'local_g1_6')
// (5, 7, 'lutff_1/in_3')
// (5, 7, 'lutff_2/in_3')
// (5, 7, 'lutff_6/in_1')
// (5, 7, 'sp4_r_v_b_2')
// (5, 7, 'sp4_r_v_b_28')
// (5, 7, 'sp4_r_v_b_6')
// (5, 8, 'sp4_r_v_b_17')
// (5, 8, 'sp4_r_v_b_39')
// (5, 9, 'local_g0_2')
// (5, 9, 'local_g1_4')
// (5, 9, 'lutff_0/in_1')
// (5, 9, 'lutff_6/in_2')
// (5, 9, 'sp4_r_v_b_26')
// (5, 9, 'sp4_r_v_b_4')
// (5, 10, 'sp4_r_v_b_15')
// (5, 10, 'sp4_r_v_b_41')
// (5, 11, 'local_g0_4')
// (5, 11, 'lutff_1/in_1')
// (5, 11, 'sp4_r_v_b_2')
// (5, 11, 'sp4_r_v_b_28')
// (5, 12, 'neigh_op_tnr_0')
// (5, 12, 'sp4_r_v_b_17')
// (5, 13, 'neigh_op_rgt_0')
// (5, 13, 'sp4_r_v_b_4')
// (5, 14, 'neigh_op_bnr_0')
// (6, 1, 'sp12_v_t_23')
// (6, 2, 'sp12_v_b_23')
// (6, 3, 'sp12_v_b_20')
// (6, 3, 'sp4_v_t_39')
// (6, 3, 'sp4_v_t_43')
// (6, 4, 'sp12_v_b_19')
// (6, 4, 'sp4_v_b_39')
// (6, 4, 'sp4_v_b_43')
// (6, 5, 'sp12_v_b_16')
// (6, 5, 'sp4_v_b_26')
// (6, 5, 'sp4_v_b_30')
// (6, 5, 'sp4_v_t_41')
// (6, 6, 'sp12_v_b_15')
// (6, 6, 'sp4_v_b_15')
// (6, 6, 'sp4_v_b_19')
// (6, 6, 'sp4_v_b_41')
// (6, 7, 'sp12_v_b_12')
// (6, 7, 'sp4_v_b_2')
// (6, 7, 'sp4_v_b_28')
// (6, 7, 'sp4_v_b_6')
// (6, 7, 'sp4_v_t_39')
// (6, 8, 'sp12_v_b_11')
// (6, 8, 'sp4_v_b_17')
// (6, 8, 'sp4_v_b_39')
// (6, 9, 'sp12_v_b_8')
// (6, 9, 'sp4_h_r_9')
// (6, 9, 'sp4_v_b_26')
// (6, 9, 'sp4_v_b_4')
// (6, 9, 'sp4_v_t_41')
// (6, 10, 'sp12_v_b_7')
// (6, 10, 'sp4_v_b_15')
// (6, 10, 'sp4_v_b_41')
// (6, 11, 'sp12_v_b_4')
// (6, 11, 'sp4_v_b_2')
// (6, 11, 'sp4_v_b_28')
// (6, 12, 'neigh_op_top_0')
// (6, 12, 'sp12_v_b_3')
// (6, 12, 'sp4_v_b_17')
// (6, 13, 'lutff_0/out')
// (6, 13, 'sp12_v_b_0')
// (6, 13, 'sp4_v_b_4')
// (6, 14, 'neigh_op_bot_0')
// (7, 9, 'local_g0_4')
// (7, 9, 'lutff_3/in_3')
// (7, 9, 'sp4_h_r_20')
// (7, 12, 'neigh_op_tnl_0')
// (7, 13, 'neigh_op_lft_0')
// (7, 14, 'neigh_op_bnl_0')
// (8, 9, 'sp4_h_r_33')
// (9, 9, 'sp4_h_r_44')
// (10, 9, 'sp4_h_l_44')

reg n264 = 0;
// (5, 5, 'neigh_op_tnr_6')
// (5, 6, 'neigh_op_rgt_6')
// (5, 7, 'neigh_op_bnr_6')
// (6, 5, 'neigh_op_top_6')
// (6, 6, 'local_g0_6')
// (6, 6, 'lutff_3/in_1')
// (6, 6, 'lutff_6/out')
// (6, 7, 'neigh_op_bot_6')
// (7, 5, 'neigh_op_tnl_6')
// (7, 6, 'neigh_op_lft_6')
// (7, 7, 'neigh_op_bnl_6')

reg n265 = 0;
// (5, 5, 'sp4_r_v_b_45')
// (5, 6, 'sp4_r_v_b_32')
// (5, 7, 'neigh_op_tnr_4')
// (5, 7, 'sp4_r_v_b_21')
// (5, 8, 'neigh_op_rgt_4')
// (5, 8, 'sp4_r_v_b_8')
// (5, 9, 'neigh_op_bnr_4')
// (6, 4, 'sp4_v_t_45')
// (6, 5, 'local_g3_5')
// (6, 5, 'lutff_1/in_3')
// (6, 5, 'sp4_v_b_45')
// (6, 6, 'sp4_v_b_32')
// (6, 7, 'neigh_op_top_4')
// (6, 7, 'sp4_v_b_21')
// (6, 8, 'lutff_4/out')
// (6, 8, 'sp4_v_b_8')
// (6, 9, 'neigh_op_bot_4')
// (7, 7, 'neigh_op_tnl_4')
// (7, 8, 'neigh_op_lft_4')
// (7, 9, 'neigh_op_bnl_4')

wire n266;
// (5, 6, 'neigh_op_tnr_1')
// (5, 7, 'neigh_op_rgt_1')
// (5, 8, 'local_g0_1')
// (5, 8, 'local_g1_1')
// (5, 8, 'lutff_0/in_2')
// (5, 8, 'lutff_2/in_2')
// (5, 8, 'lutff_3/in_2')
// (5, 8, 'lutff_6/in_2')
// (5, 8, 'neigh_op_bnr_1')
// (6, 6, 'neigh_op_top_1')
// (6, 7, 'lutff_1/out')
// (6, 8, 'neigh_op_bot_1')
// (7, 6, 'neigh_op_tnl_1')
// (7, 7, 'neigh_op_lft_1')
// (7, 8, 'neigh_op_bnl_1')

wire n267;
// (5, 6, 'neigh_op_tnr_3')
// (5, 7, 'neigh_op_rgt_3')
// (5, 8, 'neigh_op_bnr_3')
// (6, 6, 'neigh_op_top_3')
// (6, 7, 'local_g1_3')
// (6, 7, 'lutff_3/out')
// (6, 7, 'lutff_5/in_3')
// (6, 8, 'neigh_op_bot_3')
// (7, 6, 'neigh_op_tnl_3')
// (7, 7, 'neigh_op_lft_3')
// (7, 8, 'neigh_op_bnl_3')

wire n268;
// (5, 6, 'neigh_op_tnr_4')
// (5, 7, 'local_g3_4')
// (5, 7, 'lutff_1/in_0')
// (5, 7, 'neigh_op_rgt_4')
// (5, 8, 'neigh_op_bnr_4')
// (6, 6, 'neigh_op_top_4')
// (6, 7, 'local_g1_4')
// (6, 7, 'lutff_4/out')
// (6, 7, 'lutff_5/in_0')
// (6, 8, 'neigh_op_bot_4')
// (7, 6, 'neigh_op_tnl_4')
// (7, 7, 'neigh_op_lft_4')
// (7, 8, 'neigh_op_bnl_4')

wire n269;
// (5, 6, 'neigh_op_tnr_5')
// (5, 7, 'neigh_op_rgt_5')
// (5, 8, 'neigh_op_bnr_5')
// (6, 6, 'neigh_op_top_5')
// (6, 7, 'lutff_5/out')
// (6, 8, 'local_g1_5')
// (6, 8, 'lutff_0/in_2')
// (6, 8, 'lutff_3/in_3')
// (6, 8, 'neigh_op_bot_5')
// (7, 6, 'neigh_op_tnl_5')
// (7, 7, 'neigh_op_lft_5')
// (7, 8, 'neigh_op_bnl_5')

wire n270;
// (5, 6, 'neigh_op_tnr_6')
// (5, 7, 'neigh_op_rgt_6')
// (5, 8, 'local_g0_6')
// (5, 8, 'lutff_0/in_0')
// (5, 8, 'lutff_3/in_1')
// (5, 8, 'neigh_op_bnr_6')
// (6, 6, 'neigh_op_top_6')
// (6, 7, 'lutff_6/out')
// (6, 8, 'neigh_op_bot_6')
// (7, 6, 'neigh_op_tnl_6')
// (7, 7, 'neigh_op_lft_6')
// (7, 8, 'neigh_op_bnl_6')

wire n271;
// (5, 7, 'neigh_op_tnr_0')
// (5, 8, 'neigh_op_rgt_0')
// (5, 9, 'neigh_op_bnr_0')
// (6, 4, 'sp12_v_t_23')
// (6, 5, 'sp12_v_b_23')
// (6, 5, 'sp4_r_v_b_36')
// (6, 6, 'sp12_v_b_20')
// (6, 6, 'sp4_r_v_b_25')
// (6, 7, 'neigh_op_top_0')
// (6, 7, 'sp12_v_b_19')
// (6, 7, 'sp4_r_v_b_12')
// (6, 8, 'lutff_0/out')
// (6, 8, 'sp12_v_b_16')
// (6, 8, 'sp4_r_v_b_1')
// (6, 9, 'neigh_op_bot_0')
// (6, 9, 'sp12_v_b_15')
// (6, 10, 'sp12_v_b_12')
// (6, 11, 'local_g2_3')
// (6, 11, 'local_g3_3')
// (6, 11, 'lutff_2/in_3')
// (6, 11, 'lutff_6/in_3')
// (6, 11, 'lutff_7/in_3')
// (6, 11, 'sp12_v_b_11')
// (6, 12, 'sp12_v_b_8')
// (6, 13, 'sp12_v_b_7')
// (6, 14, 'sp12_v_b_4')
// (6, 15, 'sp12_v_b_3')
// (6, 16, 'sp12_v_b_0')
// (7, 4, 'sp4_v_t_36')
// (7, 5, 'sp4_v_b_36')
// (7, 6, 'sp4_v_b_25')
// (7, 7, 'neigh_op_tnl_0')
// (7, 7, 'sp4_v_b_12')
// (7, 8, 'local_g0_0')
// (7, 8, 'lutff_4/in_2')
// (7, 8, 'neigh_op_lft_0')
// (7, 8, 'sp4_h_r_7')
// (7, 8, 'sp4_v_b_1')
// (7, 9, 'neigh_op_bnl_0')
// (8, 8, 'sp4_h_r_18')
// (9, 8, 'sp4_h_r_31')
// (10, 8, 'sp4_h_r_42')
// (10, 9, 'sp4_r_v_b_42')
// (10, 10, 'sp4_r_v_b_31')
// (10, 11, 'sp4_r_v_b_18')
// (10, 12, 'sp4_r_v_b_7')
// (11, 8, 'sp4_h_l_42')
// (11, 8, 'sp4_v_t_42')
// (11, 9, 'sp4_v_b_42')
// (11, 10, 'sp4_v_b_31')
// (11, 11, 'local_g0_2')
// (11, 11, 'lutff_7/in_3')
// (11, 11, 'sp4_v_b_18')
// (11, 12, 'sp4_v_b_7')

reg n272 = 0;
// (5, 7, 'neigh_op_tnr_6')
// (5, 8, 'neigh_op_rgt_6')
// (5, 9, 'neigh_op_bnr_6')
// (6, 7, 'neigh_op_top_6')
// (6, 8, 'local_g1_6')
// (6, 8, 'lutff_6/out')
// (6, 8, 'lutff_7/in_0')
// (6, 9, 'neigh_op_bot_6')
// (7, 7, 'neigh_op_tnl_6')
// (7, 8, 'neigh_op_lft_6')
// (7, 9, 'neigh_op_bnl_6')

reg n273 = 0;
// (5, 7, 'neigh_op_tnr_7')
// (5, 8, 'neigh_op_rgt_7')
// (5, 9, 'neigh_op_bnr_7')
// (6, 7, 'neigh_op_top_7')
// (6, 8, 'local_g0_7')
// (6, 8, 'lutff_5/in_0')
// (6, 8, 'lutff_7/out')
// (6, 9, 'neigh_op_bot_7')
// (7, 7, 'neigh_op_tnl_7')
// (7, 8, 'neigh_op_lft_7')
// (7, 9, 'neigh_op_bnl_7')

wire n274;
// (5, 8, 'neigh_op_tnr_1')
// (5, 9, 'neigh_op_rgt_1')
// (5, 10, 'neigh_op_bnr_1')
// (6, 8, 'neigh_op_top_1')
// (6, 9, 'lutff_1/out')
// (6, 10, 'neigh_op_bot_1')
// (7, 8, 'neigh_op_tnl_1')
// (7, 9, 'local_g1_1')
// (7, 9, 'lutff_1/in_1')
// (7, 9, 'lutff_7/in_1')
// (7, 9, 'neigh_op_lft_1')
// (7, 10, 'neigh_op_bnl_1')

reg n275 = 0;
// (5, 8, 'neigh_op_tnr_2')
// (5, 9, 'neigh_op_rgt_2')
// (5, 10, 'neigh_op_bnr_2')
// (6, 6, 'sp4_r_v_b_40')
// (6, 7, 'sp4_r_v_b_29')
// (6, 8, 'neigh_op_top_2')
// (6, 8, 'sp4_r_v_b_16')
// (6, 9, 'local_g1_2')
// (6, 9, 'local_g1_5')
// (6, 9, 'lutff_2/out')
// (6, 9, 'lutff_4/in_1')
// (6, 9, 'lutff_6/in_2')
// (6, 9, 'sp4_r_v_b_5')
// (6, 10, 'neigh_op_bot_2')
// (7, 5, 'sp4_v_t_40')
// (7, 6, 'sp4_v_b_40')
// (7, 7, 'sp4_v_b_29')
// (7, 8, 'neigh_op_tnl_2')
// (7, 8, 'sp4_v_b_16')
// (7, 9, 'neigh_op_lft_2')
// (7, 9, 'sp4_v_b_5')
// (7, 10, 'neigh_op_bnl_2')

reg n276 = 0;
// (5, 8, 'neigh_op_tnr_3')
// (5, 9, 'neigh_op_rgt_3')
// (5, 10, 'neigh_op_bnr_3')
// (6, 8, 'neigh_op_top_3')
// (6, 9, 'local_g1_3')
// (6, 9, 'lutff_1/in_1')
// (6, 9, 'lutff_3/out')
// (6, 10, 'neigh_op_bot_3')
// (7, 8, 'neigh_op_tnl_3')
// (7, 9, 'neigh_op_lft_3')
// (7, 10, 'neigh_op_bnl_3')

reg n277 = 0;
// (5, 8, 'neigh_op_tnr_4')
// (5, 9, 'neigh_op_rgt_4')
// (5, 10, 'neigh_op_bnr_4')
// (6, 8, 'neigh_op_top_4')
// (6, 9, 'local_g0_4')
// (6, 9, 'local_g1_4')
// (6, 9, 'lutff_3/in_2')
// (6, 9, 'lutff_4/out')
// (6, 9, 'lutff_7/in_1')
// (6, 10, 'neigh_op_bot_4')
// (7, 8, 'neigh_op_tnl_4')
// (7, 9, 'neigh_op_lft_4')
// (7, 10, 'neigh_op_bnl_4')

reg n278 = 0;
// (5, 8, 'neigh_op_tnr_5')
// (5, 9, 'local_g2_5')
// (5, 9, 'local_g3_5')
// (5, 9, 'lutff_5/in_1')
// (5, 9, 'lutff_7/in_0')
// (5, 9, 'neigh_op_rgt_5')
// (5, 10, 'neigh_op_bnr_5')
// (6, 8, 'neigh_op_top_5')
// (6, 9, 'lutff_5/out')
// (6, 10, 'neigh_op_bot_5')
// (7, 8, 'neigh_op_tnl_5')
// (7, 9, 'neigh_op_lft_5')
// (7, 10, 'neigh_op_bnl_5')

reg n279 = 0;
// (5, 8, 'neigh_op_tnr_6')
// (5, 9, 'neigh_op_rgt_6')
// (5, 10, 'neigh_op_bnr_6')
// (6, 8, 'neigh_op_top_6')
// (6, 9, 'local_g2_6')
// (6, 9, 'lutff_3/in_1')
// (6, 9, 'lutff_6/out')
// (6, 10, 'neigh_op_bot_6')
// (7, 8, 'neigh_op_tnl_6')
// (7, 9, 'neigh_op_lft_6')
// (7, 10, 'neigh_op_bnl_6')

reg n280 = 0;
// (5, 8, 'neigh_op_tnr_7')
// (5, 9, 'neigh_op_rgt_7')
// (5, 10, 'neigh_op_bnr_7')
// (6, 8, 'neigh_op_top_7')
// (6, 9, 'local_g0_7')
// (6, 9, 'local_g1_7')
// (6, 9, 'lutff_1/in_2')
// (6, 9, 'lutff_5/in_1')
// (6, 9, 'lutff_7/out')
// (6, 10, 'neigh_op_bot_7')
// (7, 8, 'neigh_op_tnl_7')
// (7, 9, 'neigh_op_lft_7')
// (7, 10, 'neigh_op_bnl_7')

wire n281;
// (5, 9, 'local_g1_2')
// (5, 9, 'lutff_0/in_3')
// (5, 9, 'sp4_h_r_10')
// (6, 8, 'neigh_op_tnr_1')
// (6, 9, 'neigh_op_rgt_1')
// (6, 9, 'sp4_h_r_23')
// (6, 10, 'neigh_op_bnr_1')
// (7, 8, 'neigh_op_top_1')
// (7, 9, 'lutff_1/out')
// (7, 9, 'sp4_h_r_34')
// (7, 10, 'neigh_op_bot_1')
// (8, 8, 'neigh_op_tnl_1')
// (8, 9, 'neigh_op_lft_1')
// (8, 9, 'sp4_h_r_47')
// (8, 10, 'neigh_op_bnl_1')
// (9, 9, 'sp4_h_l_47')

wire n282;
// (5, 9, 'neigh_op_tnr_0')
// (5, 10, 'neigh_op_rgt_0')
// (5, 11, 'neigh_op_bnr_0')
// (6, 6, 'sp12_v_t_23')
// (6, 7, 'sp12_v_b_23')
// (6, 8, 'sp12_v_b_20')
// (6, 9, 'neigh_op_top_0')
// (6, 9, 'sp12_v_b_19')
// (6, 10, 'lutff_0/out')
// (6, 10, 'sp12_v_b_16')
// (6, 11, 'neigh_op_bot_0')
// (6, 11, 'sp12_v_b_15')
// (6, 12, 'sp12_v_b_12')
// (6, 13, 'local_g2_3')
// (6, 13, 'local_g3_3')
// (6, 13, 'lutff_0/in_1')
// (6, 13, 'lutff_3/in_1')
// (6, 13, 'sp12_v_b_11')
// (6, 14, 'sp12_v_b_8')
// (6, 15, 'sp12_v_b_7')
// (6, 16, 'sp12_v_b_4')
// (6, 17, 'span12_vert_3')
// (7, 9, 'neigh_op_tnl_0')
// (7, 10, 'neigh_op_lft_0')
// (7, 11, 'neigh_op_bnl_0')

reg n283 = 0;
// (5, 9, 'neigh_op_tnr_1')
// (5, 10, 'neigh_op_rgt_1')
// (5, 11, 'neigh_op_bnr_1')
// (6, 9, 'neigh_op_top_1')
// (6, 10, 'local_g0_1')
// (6, 10, 'lutff_1/out')
// (6, 10, 'lutff_4/in_1')
// (6, 10, 'lutff_5/in_2')
// (6, 11, 'neigh_op_bot_1')
// (7, 9, 'neigh_op_tnl_1')
// (7, 10, 'neigh_op_lft_1')
// (7, 11, 'neigh_op_bnl_1')

reg n284 = 0;
// (5, 9, 'neigh_op_tnr_2')
// (5, 10, 'neigh_op_rgt_2')
// (5, 11, 'neigh_op_bnr_2')
// (6, 0, 'span12_vert_23')
// (6, 1, 'sp12_v_b_23')
// (6, 2, 'sp12_v_b_20')
// (6, 3, 'sp12_v_b_19')
// (6, 4, 'sp12_v_b_16')
// (6, 5, 'sp12_v_b_15')
// (6, 6, 'sp12_v_b_12')
// (6, 7, 'sp12_v_b_11')
// (6, 8, 'local_g3_0')
// (6, 8, 'lutff_6/in_3')
// (6, 8, 'sp12_v_b_8')
// (6, 9, 'neigh_op_top_2')
// (6, 9, 'sp12_v_b_7')
// (6, 10, 'lutff_2/out')
// (6, 10, 'sp12_v_b_4')
// (6, 11, 'neigh_op_bot_2')
// (6, 11, 'sp12_v_b_3')
// (6, 12, 'sp12_v_b_0')
// (7, 9, 'neigh_op_tnl_2')
// (7, 10, 'neigh_op_lft_2')
// (7, 11, 'neigh_op_bnl_2')

reg n285 = 0;
// (5, 9, 'neigh_op_tnr_3')
// (5, 10, 'neigh_op_rgt_3')
// (5, 11, 'neigh_op_bnr_3')
// (6, 9, 'neigh_op_top_3')
// (6, 10, 'local_g1_3')
// (6, 10, 'lutff_3/out')
// (6, 10, 'lutff_5/in_1')
// (6, 11, 'neigh_op_bot_3')
// (7, 9, 'neigh_op_tnl_3')
// (7, 10, 'neigh_op_lft_3')
// (7, 11, 'neigh_op_bnl_3')

reg n286 = 0;
// (5, 9, 'neigh_op_tnr_4')
// (5, 10, 'neigh_op_rgt_4')
// (5, 11, 'neigh_op_bnr_4')
// (6, 9, 'neigh_op_top_4')
// (6, 10, 'local_g0_4')
// (6, 10, 'lutff_0/in_2')
// (6, 10, 'lutff_4/out')
// (6, 10, 'lutff_7/in_1')
// (6, 11, 'neigh_op_bot_4')
// (7, 9, 'neigh_op_tnl_4')
// (7, 10, 'neigh_op_lft_4')
// (7, 11, 'neigh_op_bnl_4')

reg n287 = 0;
// (5, 9, 'neigh_op_tnr_5')
// (5, 10, 'neigh_op_rgt_5')
// (5, 11, 'neigh_op_bnr_5')
// (6, 9, 'neigh_op_top_5')
// (6, 10, 'local_g0_5')
// (6, 10, 'lutff_0/in_1')
// (6, 10, 'lutff_5/out')
// (6, 11, 'neigh_op_bot_5')
// (7, 9, 'neigh_op_tnl_5')
// (7, 10, 'neigh_op_lft_5')
// (7, 11, 'neigh_op_bnl_5')

reg n288 = 0;
// (5, 9, 'neigh_op_tnr_6')
// (5, 10, 'neigh_op_rgt_6')
// (5, 11, 'neigh_op_bnr_6')
// (6, 9, 'neigh_op_top_6')
// (6, 10, 'local_g0_6')
// (6, 10, 'local_g1_6')
// (6, 10, 'lutff_1/in_1')
// (6, 10, 'lutff_3/in_2')
// (6, 10, 'lutff_6/out')
// (6, 11, 'neigh_op_bot_6')
// (7, 9, 'neigh_op_tnl_6')
// (7, 10, 'neigh_op_lft_6')
// (7, 11, 'neigh_op_bnl_6')

reg n289 = 0;
// (5, 9, 'neigh_op_tnr_7')
// (5, 10, 'local_g3_7')
// (5, 10, 'lutff_6/in_0')
// (5, 10, 'neigh_op_rgt_7')
// (5, 11, 'neigh_op_bnr_7')
// (6, 9, 'neigh_op_top_7')
// (6, 10, 'local_g1_7')
// (6, 10, 'lutff_6/in_2')
// (6, 10, 'lutff_7/out')
// (6, 11, 'neigh_op_bot_7')
// (7, 9, 'neigh_op_tnl_7')
// (7, 10, 'neigh_op_lft_7')
// (7, 11, 'neigh_op_bnl_7')

reg n290 = 0;
// (5, 10, 'local_g3_4')
// (5, 10, 'lutff_7/in_0')
// (5, 10, 'neigh_op_tnr_4')
// (5, 11, 'neigh_op_rgt_4')
// (5, 12, 'neigh_op_bnr_4')
// (6, 10, 'neigh_op_top_4')
// (6, 11, 'local_g0_4')
// (6, 11, 'lutff_4/out')
// (6, 11, 'lutff_7/in_1')
// (6, 12, 'neigh_op_bot_4')
// (7, 10, 'neigh_op_tnl_4')
// (7, 11, 'neigh_op_lft_4')
// (7, 12, 'neigh_op_bnl_4')

wire n291;
// (5, 10, 'neigh_op_tnr_0')
// (5, 11, 'neigh_op_rgt_0')
// (5, 12, 'neigh_op_bnr_0')
// (6, 10, 'neigh_op_top_0')
// (6, 11, 'local_g0_0')
// (6, 11, 'lutff_0/out')
// (6, 11, 'lutff_1/in_1')
// (6, 12, 'local_g0_0')
// (6, 12, 'lutff_7/in_1')
// (6, 12, 'neigh_op_bot_0')
// (7, 10, 'neigh_op_tnl_0')
// (7, 11, 'neigh_op_lft_0')
// (7, 12, 'neigh_op_bnl_0')

reg n292 = 0;
// (5, 10, 'neigh_op_tnr_2')
// (5, 11, 'neigh_op_rgt_2')
// (5, 12, 'neigh_op_bnr_2')
// (6, 10, 'neigh_op_top_2')
// (6, 11, 'local_g0_2')
// (6, 11, 'local_g1_2')
// (6, 11, 'lutff_0/in_2')
// (6, 11, 'lutff_2/out')
// (6, 11, 'lutff_4/in_1')
// (6, 12, 'neigh_op_bot_2')
// (7, 10, 'neigh_op_tnl_2')
// (7, 11, 'neigh_op_lft_2')
// (7, 12, 'neigh_op_bnl_2')

reg n293 = 0;
// (5, 10, 'neigh_op_tnr_3')
// (5, 11, 'neigh_op_rgt_3')
// (5, 12, 'neigh_op_bnr_3')
// (6, 10, 'neigh_op_top_3')
// (6, 11, 'local_g1_3')
// (6, 11, 'lutff_3/out')
// (6, 11, 'lutff_5/in_1')
// (6, 12, 'neigh_op_bot_3')
// (7, 10, 'neigh_op_tnl_3')
// (7, 11, 'neigh_op_lft_3')
// (7, 12, 'neigh_op_bnl_3')

reg n294 = 0;
// (5, 10, 'neigh_op_tnr_5')
// (5, 11, 'neigh_op_rgt_5')
// (5, 12, 'neigh_op_bnr_5')
// (6, 10, 'neigh_op_top_5')
// (6, 11, 'local_g2_5')
// (6, 11, 'lutff_0/in_1')
// (6, 11, 'lutff_5/out')
// (6, 12, 'neigh_op_bot_5')
// (7, 10, 'neigh_op_tnl_5')
// (7, 11, 'neigh_op_lft_5')
// (7, 12, 'neigh_op_bnl_5')

reg n295 = 0;
// (5, 10, 'neigh_op_tnr_6')
// (5, 11, 'neigh_op_rgt_6')
// (5, 12, 'neigh_op_bnr_6')
// (6, 10, 'neigh_op_top_6')
// (6, 11, 'local_g1_6')
// (6, 11, 'lutff_2/in_1')
// (6, 11, 'lutff_5/in_2')
// (6, 11, 'lutff_6/out')
// (6, 12, 'neigh_op_bot_6')
// (7, 10, 'neigh_op_tnl_6')
// (7, 11, 'neigh_op_lft_6')
// (7, 12, 'neigh_op_bnl_6')

reg n296 = 0;
// (5, 10, 'neigh_op_tnr_7')
// (5, 11, 'neigh_op_rgt_7')
// (5, 12, 'neigh_op_bnr_7')
// (6, 10, 'neigh_op_top_7')
// (6, 11, 'local_g0_7')
// (6, 11, 'lutff_3/in_2')
// (6, 11, 'lutff_6/in_1')
// (6, 11, 'lutff_7/out')
// (6, 12, 'neigh_op_bot_7')
// (7, 10, 'neigh_op_tnl_7')
// (7, 11, 'neigh_op_lft_7')
// (7, 12, 'neigh_op_bnl_7')

wire n297;
// (5, 11, 'neigh_op_tnr_0')
// (5, 12, 'neigh_op_rgt_0')
// (5, 13, 'neigh_op_bnr_0')
// (6, 9, 'sp4_r_v_b_36')
// (6, 10, 'sp4_r_v_b_25')
// (6, 11, 'local_g2_4')
// (6, 11, 'lutff_1/in_3')
// (6, 11, 'neigh_op_top_0')
// (6, 11, 'sp4_r_v_b_12')
// (6, 12, 'lutff_0/out')
// (6, 12, 'sp4_r_v_b_1')
// (6, 13, 'neigh_op_bot_0')
// (7, 8, 'sp4_v_t_36')
// (7, 9, 'sp4_v_b_36')
// (7, 10, 'sp4_v_b_25')
// (7, 11, 'neigh_op_tnl_0')
// (7, 11, 'sp4_v_b_12')
// (7, 12, 'neigh_op_lft_0')
// (7, 12, 'sp4_v_b_1')
// (7, 13, 'neigh_op_bnl_0')

reg n298 = 0;
// (5, 11, 'neigh_op_tnr_2')
// (5, 12, 'neigh_op_rgt_2')
// (5, 13, 'neigh_op_bnr_2')
// (6, 11, 'neigh_op_top_2')
// (6, 12, 'lutff_2/out')
// (6, 13, 'neigh_op_bot_2')
// (7, 11, 'neigh_op_tnl_2')
// (7, 12, 'local_g1_2')
// (7, 12, 'lutff_3/in_0')
// (7, 12, 'neigh_op_lft_2')
// (7, 13, 'neigh_op_bnl_2')

reg n299 = 0;
// (5, 11, 'neigh_op_tnr_3')
// (5, 12, 'neigh_op_rgt_3')
// (5, 13, 'neigh_op_bnr_3')
// (6, 11, 'neigh_op_top_3')
// (6, 12, 'local_g1_3')
// (6, 12, 'lutff_3/out')
// (6, 12, 'lutff_6/in_0')
// (6, 13, 'neigh_op_bot_3')
// (7, 11, 'neigh_op_tnl_3')
// (7, 12, 'neigh_op_lft_3')
// (7, 13, 'neigh_op_bnl_3')

reg n300 = 0;
// (5, 11, 'neigh_op_tnr_5')
// (5, 12, 'neigh_op_rgt_5')
// (5, 13, 'neigh_op_bnr_5')
// (6, 11, 'neigh_op_top_5')
// (6, 12, 'local_g0_5')
// (6, 12, 'lutff_3/in_0')
// (6, 12, 'lutff_5/out')
// (6, 13, 'neigh_op_bot_5')
// (7, 11, 'neigh_op_tnl_5')
// (7, 12, 'neigh_op_lft_5')
// (7, 13, 'neigh_op_bnl_5')

reg n301 = 0;
// (5, 11, 'neigh_op_tnr_6')
// (5, 12, 'neigh_op_rgt_6')
// (5, 13, 'neigh_op_bnr_6')
// (6, 11, 'neigh_op_top_6')
// (6, 12, 'local_g0_6')
// (6, 12, 'local_g1_6')
// (6, 12, 'lutff_1/in_1')
// (6, 12, 'lutff_2/in_1')
// (6, 12, 'lutff_6/out')
// (6, 13, 'neigh_op_bot_6')
// (7, 11, 'neigh_op_tnl_6')
// (7, 12, 'neigh_op_lft_6')
// (7, 13, 'neigh_op_bnl_6')

reg n302 = 0;
// (5, 11, 'neigh_op_tnr_7')
// (5, 12, 'neigh_op_rgt_7')
// (5, 13, 'neigh_op_bnr_7')
// (6, 11, 'neigh_op_top_7')
// (6, 12, 'local_g0_7')
// (6, 12, 'lutff_5/in_0')
// (6, 12, 'lutff_7/out')
// (6, 13, 'neigh_op_bot_7')
// (7, 11, 'neigh_op_tnl_7')
// (7, 12, 'neigh_op_lft_7')
// (7, 13, 'neigh_op_bnl_7')

reg n303 = 0;
// (5, 11, 'sp4_r_v_b_38')
// (5, 12, 'neigh_op_tnr_7')
// (5, 12, 'sp4_r_v_b_27')
// (5, 13, 'neigh_op_rgt_7')
// (5, 13, 'sp4_r_v_b_14')
// (5, 14, 'neigh_op_bnr_7')
// (5, 14, 'sp4_r_v_b_3')
// (6, 10, 'sp4_v_t_38')
// (6, 11, 'sp4_v_b_38')
// (6, 12, 'neigh_op_top_7')
// (6, 12, 'sp4_v_b_27')
// (6, 13, 'lutff_7/out')
// (6, 13, 'sp4_v_b_14')
// (6, 14, 'local_g1_3')
// (6, 14, 'lutff_5/in_1')
// (6, 14, 'neigh_op_bot_7')
// (6, 14, 'sp4_v_b_3')
// (7, 12, 'neigh_op_tnl_7')
// (7, 13, 'local_g1_7')
// (7, 13, 'lutff_4/in_0')
// (7, 13, 'neigh_op_lft_7')
// (7, 14, 'neigh_op_bnl_7')

wire n304;
// (5, 11, 'sp4_r_v_b_39')
// (5, 12, 'sp4_r_v_b_26')
// (5, 13, 'neigh_op_tnr_1')
// (5, 13, 'sp4_r_v_b_15')
// (5, 14, 'neigh_op_rgt_1')
// (5, 14, 'sp4_r_v_b_2')
// (5, 15, 'neigh_op_bnr_1')
// (6, 10, 'sp4_v_t_39')
// (6, 11, 'sp4_v_b_39')
// (6, 12, 'sp4_v_b_26')
// (6, 13, 'local_g0_7')
// (6, 13, 'lutff_0/in_3')
// (6, 13, 'neigh_op_top_1')
// (6, 13, 'sp4_v_b_15')
// (6, 14, 'lutff_1/out')
// (6, 14, 'sp4_v_b_2')
// (6, 15, 'neigh_op_bot_1')
// (7, 13, 'neigh_op_tnl_1')
// (7, 14, 'neigh_op_lft_1')
// (7, 15, 'neigh_op_bnl_1')

reg n305 = 0;
// (5, 12, 'neigh_op_tnr_1')
// (5, 13, 'neigh_op_rgt_1')
// (5, 14, 'neigh_op_bnr_1')
// (6, 12, 'neigh_op_top_1')
// (6, 13, 'local_g1_1')
// (6, 13, 'lutff_1/out')
// (6, 13, 'lutff_6/in_0')
// (6, 14, 'neigh_op_bot_1')
// (7, 12, 'neigh_op_tnl_1')
// (7, 13, 'neigh_op_lft_1')
// (7, 14, 'neigh_op_bnl_1')

reg n306 = 0;
// (5, 12, 'neigh_op_tnr_2')
// (5, 13, 'neigh_op_rgt_2')
// (5, 14, 'neigh_op_bnr_2')
// (6, 12, 'neigh_op_top_2')
// (6, 13, 'local_g1_2')
// (6, 13, 'lutff_1/in_0')
// (6, 13, 'lutff_2/out')
// (6, 14, 'neigh_op_bot_2')
// (7, 12, 'neigh_op_tnl_2')
// (7, 13, 'neigh_op_lft_2')
// (7, 14, 'neigh_op_bnl_2')

reg n307 = 0;
// (5, 12, 'neigh_op_tnr_4')
// (5, 13, 'neigh_op_rgt_4')
// (5, 14, 'neigh_op_bnr_4')
// (6, 12, 'local_g0_4')
// (6, 12, 'local_g1_4')
// (6, 12, 'lutff_0/in_0')
// (6, 12, 'lutff_2/in_0')
// (6, 12, 'lutff_7/in_0')
// (6, 12, 'neigh_op_top_4')
// (6, 13, 'local_g2_4')
// (6, 13, 'lutff_2/in_0')
// (6, 13, 'lutff_4/out')
// (6, 14, 'neigh_op_bot_4')
// (7, 12, 'neigh_op_tnl_4')
// (7, 13, 'neigh_op_lft_4')
// (7, 14, 'neigh_op_bnl_4')

reg n308 = 0;
// (5, 12, 'neigh_op_tnr_6')
// (5, 13, 'neigh_op_rgt_6')
// (5, 14, 'neigh_op_bnr_6')
// (6, 12, 'neigh_op_top_6')
// (6, 13, 'local_g0_6')
// (6, 13, 'lutff_4/in_0')
// (6, 13, 'lutff_6/out')
// (6, 14, 'neigh_op_bot_6')
// (7, 12, 'neigh_op_tnl_6')
// (7, 13, 'neigh_op_lft_6')
// (7, 14, 'neigh_op_bnl_6')

reg n309 = 0;
// (5, 12, 'sp4_r_v_b_44')
// (5, 13, 'sp4_r_v_b_33')
// (5, 14, 'sp4_r_v_b_20')
// (5, 15, 'sp4_r_v_b_9')
// (6, 6, 'sp4_h_r_7')
// (6, 11, 'local_g0_1')
// (6, 11, 'lutff_1/in_2')
// (6, 11, 'sp4_h_r_9')
// (6, 11, 'sp4_v_t_44')
// (6, 12, 'local_g3_4')
// (6, 12, 'lutff_7/in_2')
// (6, 12, 'sp4_v_b_44')
// (6, 13, 'sp4_v_b_33')
// (6, 14, 'sp4_v_b_20')
// (6, 15, 'sp4_v_b_9')
// (7, 6, 'local_g0_2')
// (7, 6, 'lutff_2/in_0')
// (7, 6, 'sp4_h_r_18')
// (7, 11, 'sp4_h_r_20')
// (8, 6, 'sp4_h_r_31')
// (8, 9, 'neigh_op_tnr_0')
// (8, 10, 'neigh_op_rgt_0')
// (8, 11, 'neigh_op_bnr_0')
// (8, 11, 'sp4_h_r_33')
// (9, 6, 'sp4_h_r_42')
// (9, 7, 'sp4_r_v_b_36')
// (9, 8, 'sp4_r_v_b_25')
// (9, 8, 'sp4_r_v_b_41')
// (9, 9, 'neigh_op_top_0')
// (9, 9, 'sp4_r_v_b_12')
// (9, 9, 'sp4_r_v_b_28')
// (9, 10, 'local_g3_0')
// (9, 10, 'lutff_0/out')
// (9, 10, 'lutff_7/in_0')
// (9, 10, 'sp4_r_v_b_1')
// (9, 10, 'sp4_r_v_b_17')
// (9, 11, 'neigh_op_bot_0')
// (9, 11, 'sp4_h_r_44')
// (9, 11, 'sp4_r_v_b_4')
// (10, 6, 'sp4_h_l_42')
// (10, 6, 'sp4_v_t_36')
// (10, 7, 'sp4_v_b_36')
// (10, 7, 'sp4_v_t_41')
// (10, 8, 'sp4_v_b_25')
// (10, 8, 'sp4_v_b_41')
// (10, 9, 'neigh_op_tnl_0')
// (10, 9, 'sp4_v_b_12')
// (10, 9, 'sp4_v_b_28')
// (10, 10, 'neigh_op_lft_0')
// (10, 10, 'sp4_v_b_1')
// (10, 10, 'sp4_v_b_17')
// (10, 11, 'neigh_op_bnl_0')
// (10, 11, 'sp4_h_l_44')
// (10, 11, 'sp4_v_b_4')

reg n310 = 0;
// (5, 12, 'sp4_r_v_b_47')
// (5, 13, 'sp4_r_v_b_34')
// (5, 14, 'neigh_op_tnr_5')
// (5, 14, 'sp4_r_v_b_23')
// (5, 15, 'neigh_op_rgt_5')
// (5, 15, 'sp4_r_v_b_10')
// (5, 16, 'neigh_op_bnr_5')
// (6, 11, 'sp4_v_t_47')
// (6, 12, 'sp4_v_b_47')
// (6, 13, 'sp4_v_b_34')
// (6, 14, 'local_g1_7')
// (6, 14, 'lutff_0/in_0')
// (6, 14, 'neigh_op_top_5')
// (6, 14, 'sp4_v_b_23')
// (6, 15, 'local_g1_5')
// (6, 15, 'lutff_5/out')
// (6, 15, 'lutff_7/in_1')
// (6, 15, 'sp4_v_b_10')
// (6, 16, 'neigh_op_bot_5')
// (7, 14, 'neigh_op_tnl_5')
// (7, 15, 'neigh_op_lft_5')
// (7, 16, 'neigh_op_bnl_5')

wire n311;
// (5, 13, 'neigh_op_tnr_0')
// (5, 14, 'neigh_op_rgt_0')
// (5, 15, 'neigh_op_bnr_0')
// (6, 13, 'neigh_op_top_0')
// (6, 14, 'local_g2_0')
// (6, 14, 'lutff_0/out')
// (6, 14, 'lutff_1/in_3')
// (6, 15, 'neigh_op_bot_0')
// (7, 13, 'neigh_op_tnl_0')
// (7, 14, 'neigh_op_lft_0')
// (7, 15, 'neigh_op_bnl_0')

reg n312 = 0;
// (5, 13, 'neigh_op_tnr_2')
// (5, 14, 'neigh_op_rgt_2')
// (5, 15, 'neigh_op_bnr_2')
// (6, 13, 'neigh_op_top_2')
// (6, 14, 'local_g1_2')
// (6, 14, 'lutff_2/out')
// (6, 14, 'lutff_5/in_0')
// (6, 14, 'sp4_r_v_b_37')
// (6, 15, 'neigh_op_bot_2')
// (6, 15, 'sp4_r_v_b_24')
// (6, 16, 'sp4_r_v_b_13')
// (7, 13, 'local_g3_2')
// (7, 13, 'lutff_5/in_0')
// (7, 13, 'lutff_7/in_0')
// (7, 13, 'neigh_op_tnl_2')
// (7, 13, 'sp4_h_r_0')
// (7, 13, 'sp4_v_t_37')
// (7, 14, 'neigh_op_lft_2')
// (7, 14, 'sp4_v_b_37')
// (7, 15, 'neigh_op_bnl_2')
// (7, 15, 'sp4_v_b_24')
// (7, 16, 'sp4_v_b_13')
// (7, 17, 'span4_vert_0')
// (8, 13, 'local_g0_5')
// (8, 13, 'lutff_1/in_0')
// (8, 13, 'sp4_h_r_13')
// (9, 13, 'sp4_h_r_24')
// (10, 13, 'sp4_h_r_37')
// (11, 13, 'sp4_h_l_37')

reg n313 = 0;
// (5, 13, 'neigh_op_tnr_3')
// (5, 14, 'neigh_op_rgt_3')
// (5, 15, 'neigh_op_bnr_3')
// (6, 13, 'neigh_op_top_3')
// (6, 14, 'local_g3_3')
// (6, 14, 'lutff_3/out')
// (6, 14, 'lutff_4/in_0')
// (6, 15, 'neigh_op_bot_3')
// (7, 13, 'neigh_op_tnl_3')
// (7, 14, 'neigh_op_lft_3')
// (7, 15, 'neigh_op_bnl_3')

reg n314 = 0;
// (5, 13, 'neigh_op_tnr_4')
// (5, 14, 'neigh_op_rgt_4')
// (5, 15, 'neigh_op_bnr_4')
// (6, 13, 'neigh_op_top_4')
// (6, 14, 'local_g0_4')
// (6, 14, 'lutff_4/out')
// (6, 14, 'lutff_6/in_0')
// (6, 15, 'neigh_op_bot_4')
// (7, 13, 'neigh_op_tnl_4')
// (7, 14, 'neigh_op_lft_4')
// (7, 15, 'neigh_op_bnl_4')

reg n315 = 0;
// (5, 13, 'neigh_op_tnr_6')
// (5, 14, 'neigh_op_rgt_6')
// (5, 15, 'neigh_op_bnr_6')
// (6, 13, 'neigh_op_top_6')
// (6, 14, 'lutff_6/out')
// (6, 15, 'local_g1_6')
// (6, 15, 'lutff_5/in_0')
// (6, 15, 'neigh_op_bot_6')
// (7, 13, 'neigh_op_tnl_6')
// (7, 14, 'neigh_op_lft_6')
// (7, 15, 'neigh_op_bnl_6')

reg n316 = 0;
// (5, 14, 'neigh_op_tnr_0')
// (5, 15, 'neigh_op_rgt_0')
// (5, 16, 'neigh_op_bnr_0')
// (6, 14, 'neigh_op_top_0')
// (6, 15, 'local_g3_0')
// (6, 15, 'lutff_0/out')
// (6, 15, 'lutff_1/in_0')
// (6, 16, 'neigh_op_bot_0')
// (7, 14, 'neigh_op_tnl_0')
// (7, 15, 'neigh_op_lft_0')
// (7, 16, 'neigh_op_bnl_0')

reg n317 = 0;
// (5, 14, 'neigh_op_tnr_1')
// (5, 15, 'neigh_op_rgt_1')
// (5, 16, 'neigh_op_bnr_1')
// (6, 14, 'neigh_op_top_1')
// (6, 15, 'local_g1_1')
// (6, 15, 'lutff_1/out')
// (6, 15, 'lutff_4/in_0')
// (6, 16, 'neigh_op_bot_1')
// (7, 14, 'neigh_op_tnl_1')
// (7, 15, 'neigh_op_lft_1')
// (7, 16, 'neigh_op_bnl_1')

reg n318 = 0;
// (5, 14, 'neigh_op_tnr_4')
// (5, 15, 'neigh_op_rgt_4')
// (5, 16, 'neigh_op_bnr_4')
// (6, 12, 'sp4_r_v_b_44')
// (6, 13, 'local_g2_1')
// (6, 13, 'lutff_3/in_0')
// (6, 13, 'sp4_r_v_b_33')
// (6, 14, 'local_g1_4')
// (6, 14, 'lutff_1/in_0')
// (6, 14, 'lutff_3/in_0')
// (6, 14, 'neigh_op_top_4')
// (6, 14, 'sp4_r_v_b_20')
// (6, 15, 'local_g1_4')
// (6, 15, 'lutff_4/out')
// (6, 15, 'lutff_7/in_0')
// (6, 15, 'sp4_r_v_b_9')
// (6, 16, 'neigh_op_bot_4')
// (7, 11, 'sp4_v_t_44')
// (7, 12, 'sp4_v_b_44')
// (7, 13, 'sp4_v_b_33')
// (7, 14, 'neigh_op_tnl_4')
// (7, 14, 'sp4_v_b_20')
// (7, 15, 'neigh_op_lft_4')
// (7, 15, 'sp4_v_b_9')
// (7, 16, 'neigh_op_bnl_4')

reg n319 = 0;
// (5, 14, 'neigh_op_tnr_7')
// (5, 15, 'neigh_op_rgt_7')
// (5, 16, 'neigh_op_bnr_7')
// (6, 14, 'neigh_op_top_7')
// (6, 15, 'local_g1_7')
// (6, 15, 'lutff_0/in_0')
// (6, 15, 'lutff_7/out')
// (6, 16, 'neigh_op_bot_7')
// (7, 14, 'neigh_op_tnl_7')
// (7, 15, 'neigh_op_lft_7')
// (7, 16, 'neigh_op_bnl_7')

wire n320;
// (6, 1, 'neigh_op_tnr_0')
// (6, 2, 'local_g2_0')
// (6, 2, 'local_g3_0')
// (6, 2, 'lutff_1/in_3')
// (6, 2, 'lutff_6/in_1')
// (6, 2, 'neigh_op_rgt_0')
// (6, 3, 'neigh_op_bnr_0')
// (7, 1, 'neigh_op_top_0')
// (7, 2, 'local_g1_0')
// (7, 2, 'lutff_0/out')
// (7, 2, 'lutff_3/in_0')
// (7, 3, 'neigh_op_bot_0')
// (8, 1, 'neigh_op_tnl_0')
// (8, 2, 'neigh_op_lft_0')
// (8, 3, 'neigh_op_bnl_0')

wire n321;
// (6, 1, 'neigh_op_tnr_1')
// (6, 2, 'neigh_op_rgt_1')
// (6, 3, 'neigh_op_bnr_1')
// (7, 1, 'neigh_op_top_1')
// (7, 2, 'local_g1_1')
// (7, 2, 'lutff_1/out')
// (7, 2, 'lutff_2/in_0')
// (7, 2, 'lutff_4/in_2')
// (7, 2, 'lutff_6/in_2')
// (7, 3, 'neigh_op_bot_1')
// (8, 1, 'neigh_op_tnl_1')
// (8, 2, 'neigh_op_lft_1')
// (8, 3, 'neigh_op_bnl_1')

wire n322;
// (6, 1, 'neigh_op_tnr_2')
// (6, 2, 'local_g2_2')
// (6, 2, 'local_g3_2')
// (6, 2, 'lutff_1/in_2')
// (6, 2, 'lutff_2/in_2')
// (6, 2, 'neigh_op_rgt_2')
// (6, 3, 'neigh_op_bnr_2')
// (7, 1, 'neigh_op_top_2')
// (7, 2, 'lutff_2/out')
// (7, 3, 'neigh_op_bot_2')
// (8, 1, 'neigh_op_tnl_2')
// (8, 2, 'neigh_op_lft_2')
// (8, 3, 'neigh_op_bnl_2')

wire n323;
// (6, 1, 'neigh_op_tnr_3')
// (6, 2, 'neigh_op_rgt_3')
// (6, 3, 'neigh_op_bnr_3')
// (7, 1, 'neigh_op_top_3')
// (7, 2, 'local_g2_3')
// (7, 2, 'lutff_2/in_1')
// (7, 2, 'lutff_3/out')
// (7, 2, 'lutff_4/in_3')
// (7, 3, 'neigh_op_bot_3')
// (8, 1, 'neigh_op_tnl_3')
// (8, 2, 'neigh_op_lft_3')
// (8, 3, 'neigh_op_bnl_3')

wire n324;
// (6, 1, 'neigh_op_tnr_4')
// (6, 2, 'neigh_op_rgt_4')
// (6, 3, 'local_g0_4')
// (6, 3, 'local_g1_4')
// (6, 3, 'lutff_0/in_3')
// (6, 3, 'lutff_1/in_2')
// (6, 3, 'lutff_2/in_1')
// (6, 3, 'lutff_3/in_0')
// (6, 3, 'lutff_5/in_3')
// (6, 3, 'lutff_6/in_1')
// (6, 3, 'lutff_7/in_2')
// (6, 3, 'neigh_op_bnr_4')
// (7, 1, 'neigh_op_top_4')
// (7, 2, 'lutff_4/out')
// (7, 3, 'neigh_op_bot_4')
// (8, 1, 'neigh_op_tnl_4')
// (8, 2, 'neigh_op_lft_4')
// (8, 3, 'neigh_op_bnl_4')

wire n325;
// (6, 1, 'neigh_op_tnr_6')
// (6, 2, 'local_g2_6')
// (6, 2, 'local_g3_6')
// (6, 2, 'lutff_1/in_1')
// (6, 2, 'lutff_2/in_1')
// (6, 2, 'neigh_op_rgt_6')
// (6, 3, 'local_g0_6')
// (6, 3, 'local_g1_6')
// (6, 3, 'lutff_0/in_2')
// (6, 3, 'lutff_1/in_3')
// (6, 3, 'lutff_2/in_0')
// (6, 3, 'lutff_3/in_1')
// (6, 3, 'lutff_5/in_0')
// (6, 3, 'lutff_6/in_0')
// (6, 3, 'lutff_7/in_3')
// (6, 3, 'neigh_op_bnr_6')
// (7, 1, 'neigh_op_top_6')
// (7, 2, 'lutff_6/out')
// (7, 3, 'neigh_op_bot_6')
// (8, 1, 'neigh_op_tnl_6')
// (8, 2, 'neigh_op_lft_6')
// (8, 3, 'neigh_op_bnl_6')

wire n326;
// (6, 1, 'neigh_op_tnr_7')
// (6, 2, 'local_g2_7')
// (6, 2, 'local_g3_7')
// (6, 2, 'lutff_3/in_0')
// (6, 2, 'lutff_5/in_1')
// (6, 2, 'neigh_op_rgt_7')
// (6, 3, 'neigh_op_bnr_7')
// (7, 1, 'neigh_op_top_7')
// (7, 2, 'lutff_7/out')
// (7, 3, 'neigh_op_bot_7')
// (8, 1, 'neigh_op_tnl_7')
// (8, 2, 'neigh_op_lft_7')
// (8, 3, 'neigh_op_bnl_7')

wire n327;
// (6, 2, 'local_g0_2')
// (6, 2, 'local_g1_2')
// (6, 2, 'lutff_3/in_2')
// (6, 2, 'lutff_5/in_3')
// (6, 2, 'sp4_h_r_10')
// (7, 1, 'neigh_op_tnr_1')
// (7, 2, 'neigh_op_rgt_1')
// (7, 2, 'sp4_h_r_23')
// (7, 3, 'neigh_op_bnr_1')
// (8, 1, 'neigh_op_top_1')
// (8, 2, 'local_g0_1')
// (8, 2, 'local_g1_1')
// (8, 2, 'lutff_1/out')
// (8, 2, 'lutff_6/in_2')
// (8, 2, 'lutff_7/in_2')
// (8, 2, 'sp4_h_r_34')
// (8, 3, 'neigh_op_bot_1')
// (9, 1, 'neigh_op_tnl_1')
// (9, 2, 'neigh_op_lft_1')
// (9, 2, 'sp4_h_r_47')
// (9, 3, 'neigh_op_bnl_1')
// (10, 2, 'sp4_h_l_47')

wire n328;
// (6, 2, 'neigh_op_tnr_0')
// (6, 3, 'neigh_op_rgt_0')
// (6, 4, 'neigh_op_bnr_0')
// (7, 2, 'neigh_op_top_0')
// (7, 3, 'local_g0_0')
// (7, 3, 'lutff_0/out')
// (7, 3, 'lutff_5/in_1')
// (7, 4, 'neigh_op_bot_0')
// (8, 2, 'neigh_op_tnl_0')
// (8, 3, 'neigh_op_lft_0')
// (8, 4, 'local_g3_0')
// (8, 4, 'lutff_0/in_3')
// (8, 4, 'neigh_op_bnl_0')

wire n329;
// (6, 2, 'neigh_op_tnr_1')
// (6, 3, 'neigh_op_rgt_1')
// (6, 4, 'neigh_op_bnr_1')
// (7, 2, 'neigh_op_top_1')
// (7, 2, 'sp4_r_v_b_46')
// (7, 3, 'lutff_1/out')
// (7, 3, 'sp4_r_v_b_35')
// (7, 4, 'local_g1_1')
// (7, 4, 'local_g3_6')
// (7, 4, 'lutff_1/in_1')
// (7, 4, 'lutff_4/in_2')
// (7, 4, 'lutff_6/in_1')
// (7, 4, 'neigh_op_bot_1')
// (7, 4, 'sp4_r_v_b_22')
// (7, 5, 'sp4_r_v_b_11')
// (8, 1, 'sp4_v_t_46')
// (8, 2, 'neigh_op_tnl_1')
// (8, 2, 'sp4_v_b_46')
// (8, 3, 'neigh_op_lft_1')
// (8, 3, 'sp4_v_b_35')
// (8, 4, 'neigh_op_bnl_1')
// (8, 4, 'sp4_v_b_22')
// (8, 5, 'sp4_v_b_11')

wire n330;
// (6, 2, 'neigh_op_tnr_2')
// (6, 3, 'neigh_op_rgt_2')
// (6, 3, 'sp4_r_v_b_36')
// (6, 4, 'neigh_op_bnr_2')
// (6, 4, 'sp4_r_v_b_25')
// (6, 5, 'sp4_r_v_b_12')
// (6, 6, 'sp4_r_v_b_1')
// (7, 2, 'neigh_op_top_2')
// (7, 2, 'sp4_v_t_36')
// (7, 3, 'lutff_2/out')
// (7, 3, 'sp4_v_b_36')
// (7, 4, 'neigh_op_bot_2')
// (7, 4, 'sp4_v_b_25')
// (7, 5, 'local_g1_4')
// (7, 5, 'lutff_3/in_2')
// (7, 5, 'sp4_v_b_12')
// (7, 6, 'sp4_v_b_1')
// (8, 2, 'neigh_op_tnl_2')
// (8, 3, 'neigh_op_lft_2')
// (8, 4, 'neigh_op_bnl_2')

wire n331;
// (6, 2, 'neigh_op_tnr_4')
// (6, 3, 'neigh_op_rgt_4')
// (6, 4, 'neigh_op_bnr_4')
// (7, 2, 'neigh_op_top_4')
// (7, 3, 'local_g0_4')
// (7, 3, 'local_g1_4')
// (7, 3, 'lutff_2/in_2')
// (7, 3, 'lutff_4/out')
// (7, 3, 'lutff_5/in_2')
// (7, 4, 'neigh_op_bot_4')
// (8, 2, 'neigh_op_tnl_4')
// (8, 3, 'neigh_op_lft_4')
// (8, 4, 'neigh_op_bnl_4')

wire n332;
// (6, 2, 'neigh_op_tnr_5')
// (6, 3, 'neigh_op_rgt_5')
// (6, 3, 'sp4_r_v_b_42')
// (6, 4, 'neigh_op_bnr_5')
// (6, 4, 'sp4_r_v_b_31')
// (6, 5, 'sp4_r_v_b_18')
// (6, 6, 'sp4_r_v_b_7')
// (7, 2, 'neigh_op_top_5')
// (7, 2, 'sp4_v_t_42')
// (7, 3, 'lutff_5/out')
// (7, 3, 'sp4_v_b_42')
// (7, 4, 'neigh_op_bot_5')
// (7, 4, 'sp4_v_b_31')
// (7, 5, 'local_g0_2')
// (7, 5, 'lutff_3/in_1')
// (7, 5, 'lutff_5/in_1')
// (7, 5, 'sp4_v_b_18')
// (7, 6, 'sp4_v_b_7')
// (8, 2, 'neigh_op_tnl_5')
// (8, 3, 'neigh_op_lft_5')
// (8, 4, 'neigh_op_bnl_5')

wire n333;
// (6, 2, 'neigh_op_tnr_6')
// (6, 3, 'neigh_op_rgt_6')
// (6, 4, 'neigh_op_bnr_6')
// (7, 2, 'neigh_op_top_6')
// (7, 3, 'lutff_6/out')
// (7, 4, 'local_g0_6')
// (7, 4, 'local_g1_6')
// (7, 4, 'lutff_1/in_3')
// (7, 4, 'lutff_2/in_3')
// (7, 4, 'neigh_op_bot_6')
// (8, 2, 'neigh_op_tnl_6')
// (8, 3, 'neigh_op_lft_6')
// (8, 4, 'neigh_op_bnl_6')

wire n334;
// (6, 2, 'neigh_op_tnr_7')
// (6, 3, 'neigh_op_rgt_7')
// (6, 4, 'neigh_op_bnr_7')
// (7, 2, 'neigh_op_top_7')
// (7, 3, 'lutff_7/out')
// (7, 4, 'local_g0_7')
// (7, 4, 'local_g1_7')
// (7, 4, 'lutff_1/in_2')
// (7, 4, 'lutff_2/in_0')
// (7, 4, 'neigh_op_bot_7')
// (8, 2, 'neigh_op_tnl_7')
// (8, 3, 'local_g1_7')
// (8, 3, 'lutff_4/in_2')
// (8, 3, 'neigh_op_lft_7')
// (8, 4, 'neigh_op_bnl_7')

wire n335;
// (6, 2, 'sp4_h_r_6')
// (7, 1, 'neigh_op_tnr_7')
// (7, 2, 'local_g0_3')
// (7, 2, 'local_g1_3')
// (7, 2, 'lutff_2/in_2')
// (7, 2, 'lutff_6/in_3')
// (7, 2, 'neigh_op_rgt_7')
// (7, 2, 'sp4_h_r_19')
// (7, 3, 'neigh_op_bnr_7')
// (8, 1, 'neigh_op_top_7')
// (8, 2, 'lutff_7/out')
// (8, 2, 'sp4_h_r_30')
// (8, 3, 'neigh_op_bot_7')
// (9, 1, 'neigh_op_tnl_7')
// (9, 2, 'neigh_op_lft_7')
// (9, 2, 'sp4_h_r_43')
// (9, 3, 'neigh_op_bnl_7')
// (10, 2, 'sp4_h_l_43')

wire n336;
// (6, 2, 'sp4_r_v_b_44')
// (6, 3, 'neigh_op_tnr_2')
// (6, 3, 'sp4_r_v_b_33')
// (6, 4, 'neigh_op_rgt_2')
// (6, 4, 'sp4_r_v_b_20')
// (6, 5, 'neigh_op_bnr_2')
// (6, 5, 'sp4_r_v_b_9')
// (7, 1, 'sp4_v_t_44')
// (7, 2, 'sp4_v_b_44')
// (7, 3, 'neigh_op_top_2')
// (7, 3, 'sp4_v_b_33')
// (7, 4, 'local_g0_2')
// (7, 4, 'lutff_2/out')
// (7, 4, 'lutff_4/in_0')
// (7, 4, 'lutff_6/in_0')
// (7, 4, 'sp4_v_b_20')
// (7, 5, 'local_g1_1')
// (7, 5, 'local_g1_2')
// (7, 5, 'lutff_2/in_1')
// (7, 5, 'lutff_3/in_3')
// (7, 5, 'neigh_op_bot_2')
// (7, 5, 'sp4_v_b_9')
// (8, 3, 'neigh_op_tnl_2')
// (8, 4, 'neigh_op_lft_2')
// (8, 5, 'neigh_op_bnl_2')

wire n337;
// (6, 3, 'neigh_op_tnr_0')
// (6, 4, 'local_g2_0')
// (6, 4, 'local_g3_0')
// (6, 4, 'lutff_1/in_3')
// (6, 4, 'lutff_7/in_2')
// (6, 4, 'neigh_op_rgt_0')
// (6, 5, 'neigh_op_bnr_0')
// (7, 3, 'neigh_op_top_0')
// (7, 4, 'local_g1_0')
// (7, 4, 'lutff_0/out')
// (7, 4, 'lutff_3/in_0')
// (7, 5, 'neigh_op_bot_0')
// (8, 3, 'neigh_op_tnl_0')
// (8, 4, 'neigh_op_lft_0')
// (8, 5, 'neigh_op_bnl_0')

wire n338;
// (6, 3, 'neigh_op_tnr_1')
// (6, 4, 'neigh_op_rgt_1')
// (6, 5, 'local_g1_1')
// (6, 5, 'lutff_1/in_1')
// (6, 5, 'neigh_op_bnr_1')
// (7, 3, 'neigh_op_top_1')
// (7, 4, 'lutff_1/out')
// (7, 5, 'neigh_op_bot_1')
// (8, 3, 'neigh_op_tnl_1')
// (8, 4, 'neigh_op_lft_1')
// (8, 5, 'neigh_op_bnl_1')

wire n339;
// (6, 3, 'neigh_op_tnr_4')
// (6, 4, 'neigh_op_rgt_4')
// (6, 5, 'neigh_op_bnr_4')
// (7, 1, 'sp4_r_v_b_44')
// (7, 2, 'sp4_r_v_b_33')
// (7, 3, 'neigh_op_top_4')
// (7, 3, 'sp4_r_v_b_20')
// (7, 4, 'lutff_4/out')
// (7, 4, 'sp4_r_v_b_9')
// (7, 5, 'neigh_op_bot_4')
// (7, 5, 'sp4_r_v_b_37')
// (7, 6, 'sp4_r_v_b_24')
// (7, 7, 'sp4_r_v_b_13')
// (7, 8, 'sp4_r_v_b_0')
// (8, 0, 'span4_vert_44')
// (8, 1, 'sp4_v_b_44')
// (8, 2, 'sp4_v_b_33')
// (8, 3, 'neigh_op_tnl_4')
// (8, 3, 'sp4_v_b_20')
// (8, 4, 'neigh_op_lft_4')
// (8, 4, 'sp4_v_b_9')
// (8, 4, 'sp4_v_t_37')
// (8, 5, 'neigh_op_bnl_4')
// (8, 5, 'sp4_v_b_37')
// (8, 6, 'sp4_v_b_24')
// (8, 7, 'sp4_v_b_13')
// (8, 8, 'local_g0_0')
// (8, 8, 'lutff_0/in_2')
// (8, 8, 'sp4_v_b_0')

wire n340;
// (6, 3, 'neigh_op_tnr_5')
// (6, 4, 'neigh_op_rgt_5')
// (6, 5, 'neigh_op_bnr_5')
// (7, 3, 'neigh_op_top_5')
// (7, 4, 'local_g0_5')
// (7, 4, 'local_g1_5')
// (7, 4, 'lutff_2/in_2')
// (7, 4, 'lutff_3/in_2')
// (7, 4, 'lutff_5/out')
// (7, 5, 'neigh_op_bot_5')
// (8, 3, 'neigh_op_tnl_5')
// (8, 4, 'neigh_op_lft_5')
// (8, 5, 'neigh_op_bnl_5')

wire n341;
// (6, 3, 'neigh_op_tnr_6')
// (6, 4, 'neigh_op_rgt_6')
// (6, 4, 'sp4_r_v_b_44')
// (6, 5, 'neigh_op_bnr_6')
// (6, 5, 'sp4_r_v_b_33')
// (6, 6, 'sp4_r_v_b_20')
// (6, 7, 'sp4_r_v_b_9')
// (7, 3, 'neigh_op_top_6')
// (7, 3, 'sp4_v_t_44')
// (7, 4, 'lutff_6/out')
// (7, 4, 'sp4_v_b_44')
// (7, 5, 'neigh_op_bot_6')
// (7, 5, 'sp4_v_b_33')
// (7, 6, 'sp4_v_b_20')
// (7, 7, 'local_g1_1')
// (7, 7, 'lutff_0/in_2')
// (7, 7, 'sp4_v_b_9')
// (8, 3, 'neigh_op_tnl_6')
// (8, 4, 'neigh_op_lft_6')
// (8, 5, 'neigh_op_bnl_6')

wire n342;
// (6, 3, 'sp12_h_r_1')
// (7, 3, 'sp12_h_r_2')
// (8, 2, 'neigh_op_tnr_7')
// (8, 3, 'local_g2_7')
// (8, 3, 'local_g3_7')
// (8, 3, 'lutff_0/in_1')
// (8, 3, 'lutff_4/in_0')
// (8, 3, 'lutff_6/in_1')
// (8, 3, 'neigh_op_rgt_7')
// (8, 3, 'sp12_h_r_5')
// (8, 4, 'neigh_op_bnr_7')
// (9, 2, 'neigh_op_top_7')
// (9, 3, 'lutff_7/out')
// (9, 3, 'sp12_h_r_6')
// (9, 4, 'neigh_op_bot_7')
// (10, 2, 'neigh_op_tnl_7')
// (10, 3, 'neigh_op_lft_7')
// (10, 3, 'sp12_h_r_9')
// (10, 4, 'neigh_op_bnl_7')
// (11, 3, 'local_g1_2')
// (11, 3, 'lutff_5/in_2')
// (11, 3, 'sp12_h_r_10')
// (12, 3, 'sp12_h_r_13')
// (13, 3, 'span12_horz_13')

wire n343;
// (6, 4, 'neigh_op_tnr_0')
// (6, 5, 'neigh_op_rgt_0')
// (6, 6, 'neigh_op_bnr_0')
// (7, 4, 'neigh_op_top_0')
// (7, 5, 'lutff_0/out')
// (7, 6, 'neigh_op_bot_0')
// (8, 4, 'neigh_op_tnl_0')
// (8, 5, 'local_g0_0')
// (8, 5, 'lutff_0/in_2')
// (8, 5, 'neigh_op_lft_0')
// (8, 6, 'neigh_op_bnl_0')

wire n344;
// (6, 4, 'neigh_op_tnr_3')
// (6, 5, 'neigh_op_rgt_3')
// (6, 6, 'neigh_op_bnr_3')
// (7, 4, 'neigh_op_top_3')
// (7, 5, 'lutff_3/out')
// (7, 6, 'neigh_op_bot_3')
// (8, 4, 'neigh_op_tnl_3')
// (8, 5, 'local_g0_3')
// (8, 5, 'lutff_0/in_1')
// (8, 5, 'neigh_op_lft_3')
// (8, 6, 'neigh_op_bnl_3')

wire n345;
// (6, 4, 'neigh_op_tnr_4')
// (6, 5, 'neigh_op_rgt_4')
// (6, 6, 'neigh_op_bnr_4')
// (7, 4, 'neigh_op_top_4')
// (7, 5, 'lutff_4/out')
// (7, 6, 'neigh_op_bot_4')
// (8, 4, 'local_g2_4')
// (8, 4, 'lutff_2/in_0')
// (8, 4, 'lutff_6/in_2')
// (8, 4, 'neigh_op_tnl_4')
// (8, 5, 'neigh_op_lft_4')
// (8, 6, 'neigh_op_bnl_4')

wire n346;
// (6, 4, 'neigh_op_tnr_5')
// (6, 5, 'neigh_op_rgt_5')
// (6, 6, 'local_g0_5')
// (6, 6, 'local_g1_5')
// (6, 6, 'lutff_3/in_2')
// (6, 6, 'lutff_6/in_2')
// (6, 6, 'neigh_op_bnr_5')
// (7, 4, 'neigh_op_top_5')
// (7, 5, 'lutff_5/out')
// (7, 6, 'neigh_op_bot_5')
// (8, 4, 'neigh_op_tnl_5')
// (8, 5, 'local_g0_5')
// (8, 5, 'lutff_7/in_0')
// (8, 5, 'neigh_op_lft_5')
// (8, 6, 'local_g2_5')
// (8, 6, 'lutff_3/in_2')
// (8, 6, 'neigh_op_bnl_5')

reg n347 = 0;
// (6, 4, 'neigh_op_tnr_6')
// (6, 5, 'neigh_op_rgt_6')
// (6, 5, 'sp4_r_v_b_44')
// (6, 6, 'neigh_op_bnr_6')
// (6, 6, 'sp4_r_v_b_33')
// (6, 7, 'sp4_r_v_b_20')
// (6, 8, 'sp4_r_v_b_9')
// (6, 9, 'sp4_r_v_b_37')
// (6, 10, 'sp4_r_v_b_24')
// (6, 11, 'sp4_r_v_b_13')
// (6, 12, 'sp4_r_v_b_0')
// (6, 13, 'sp4_r_v_b_37')
// (6, 14, 'sp4_r_v_b_24')
// (6, 15, 'sp4_r_v_b_13')
// (6, 16, 'sp4_r_v_b_0')
// (7, 4, 'neigh_op_top_6')
// (7, 4, 'sp4_v_t_44')
// (7, 5, 'lutff_6/out')
// (7, 5, 'sp4_v_b_44')
// (7, 6, 'local_g1_6')
// (7, 6, 'lutff_7/in_0')
// (7, 6, 'neigh_op_bot_6')
// (7, 6, 'sp4_v_b_33')
// (7, 7, 'sp4_v_b_20')
// (7, 8, 'sp4_v_b_9')
// (7, 8, 'sp4_v_t_37')
// (7, 9, 'sp4_v_b_37')
// (7, 10, 'sp4_v_b_24')
// (7, 11, 'local_g0_5')
// (7, 11, 'lutff_5/in_0')
// (7, 11, 'sp4_v_b_13')
// (7, 12, 'sp4_v_b_0')
// (7, 12, 'sp4_v_t_37')
// (7, 13, 'local_g2_5')
// (7, 13, 'lutff_1/in_2')
// (7, 13, 'lutff_7/in_2')
// (7, 13, 'sp4_v_b_37')
// (7, 14, 'sp4_v_b_24')
// (7, 15, 'sp4_v_b_13')
// (7, 16, 'sp4_v_b_0')
// (8, 4, 'neigh_op_tnl_6')
// (8, 5, 'neigh_op_lft_6')
// (8, 6, 'neigh_op_bnl_6')

reg n348 = 0;
// (6, 4, 'neigh_op_tnr_7')
// (6, 5, 'neigh_op_rgt_7')
// (6, 6, 'neigh_op_bnr_7')
// (7, 4, 'neigh_op_top_7')
// (7, 5, 'local_g0_7')
// (7, 5, 'lutff_2/in_3')
// (7, 5, 'lutff_7/out')
// (7, 6, 'neigh_op_bot_7')
// (8, 4, 'neigh_op_tnl_7')
// (8, 5, 'neigh_op_lft_7')
// (8, 6, 'neigh_op_bnl_7')

reg n349 = 0;
// (6, 5, 'neigh_op_tnr_2')
// (6, 6, 'neigh_op_rgt_2')
// (6, 7, 'neigh_op_bnr_2')
// (7, 5, 'neigh_op_top_2')
// (7, 6, 'lutff_2/out')
// (7, 7, 'neigh_op_bot_2')
// (8, 5, 'local_g3_2')
// (8, 5, 'lutff_6/in_3')
// (8, 5, 'neigh_op_tnl_2')
// (8, 6, 'neigh_op_lft_2')
// (8, 7, 'neigh_op_bnl_2')

reg n350 = 0;
// (6, 5, 'neigh_op_tnr_6')
// (6, 6, 'neigh_op_rgt_6')
// (6, 7, 'neigh_op_bnr_6')
// (7, 5, 'neigh_op_top_6')
// (7, 6, 'lutff_6/out')
// (7, 6, 'sp4_r_v_b_45')
// (7, 7, 'neigh_op_bot_6')
// (7, 7, 'sp4_r_v_b_32')
// (7, 8, 'sp4_r_v_b_21')
// (7, 9, 'sp4_r_v_b_8')
// (8, 5, 'neigh_op_tnl_6')
// (8, 5, 'sp4_h_r_8')
// (8, 5, 'sp4_v_t_45')
// (8, 6, 'neigh_op_lft_6')
// (8, 6, 'sp4_v_b_45')
// (8, 7, 'neigh_op_bnl_6')
// (8, 7, 'sp4_v_b_32')
// (8, 8, 'sp4_v_b_21')
// (8, 9, 'sp4_v_b_8')
// (9, 5, 'sp4_h_r_21')
// (10, 5, 'sp4_h_r_32')
// (11, 5, 'local_g2_5')
// (11, 5, 'lutff_0/in_3')
// (11, 5, 'sp4_h_r_45')
// (12, 5, 'sp4_h_l_45')

reg n351 = 0;
// (6, 5, 'neigh_op_tnr_7')
// (6, 6, 'neigh_op_rgt_7')
// (6, 7, 'neigh_op_bnr_7')
// (7, 1, 'sp12_v_t_22')
// (7, 2, 'sp12_v_b_22')
// (7, 3, 'sp12_v_b_21')
// (7, 4, 'local_g2_2')
// (7, 4, 'lutff_7/in_3')
// (7, 4, 'sp12_v_b_18')
// (7, 5, 'neigh_op_top_7')
// (7, 5, 'sp12_v_b_17')
// (7, 6, 'lutff_7/out')
// (7, 6, 'sp12_v_b_14')
// (7, 7, 'neigh_op_bot_7')
// (7, 7, 'sp12_v_b_13')
// (7, 8, 'sp12_v_b_10')
// (7, 9, 'sp12_v_b_9')
// (7, 10, 'sp12_v_b_6')
// (7, 11, 'sp12_v_b_5')
// (7, 12, 'sp12_v_b_2')
// (7, 13, 'sp12_v_b_1')
// (8, 5, 'neigh_op_tnl_7')
// (8, 6, 'neigh_op_lft_7')
// (8, 7, 'neigh_op_bnl_7')

reg n352 = 0;
// (6, 6, 'neigh_op_tnr_5')
// (6, 7, 'neigh_op_rgt_5')
// (6, 8, 'neigh_op_bnr_5')
// (7, 6, 'neigh_op_top_5')
// (7, 7, 'local_g0_5')
// (7, 7, 'lutff_5/out')
// (7, 7, 'lutff_7/in_0')
// (7, 8, 'neigh_op_bot_5')
// (8, 6, 'neigh_op_tnl_5')
// (8, 7, 'neigh_op_lft_5')
// (8, 8, 'neigh_op_bnl_5')

reg n353 = 0;
// (6, 6, 'neigh_op_tnr_7')
// (6, 7, 'neigh_op_rgt_7')
// (6, 8, 'neigh_op_bnr_7')
// (7, 5, 'local_g2_7')
// (7, 5, 'lutff_4/in_3')
// (7, 5, 'sp4_r_v_b_39')
// (7, 6, 'neigh_op_top_7')
// (7, 6, 'sp4_r_v_b_26')
// (7, 7, 'local_g0_7')
// (7, 7, 'lutff_3/in_0')
// (7, 7, 'lutff_7/out')
// (7, 7, 'sp4_r_v_b_15')
// (7, 8, 'neigh_op_bot_7')
// (7, 8, 'sp4_r_v_b_2')
// (8, 4, 'sp4_v_t_39')
// (8, 5, 'sp4_v_b_39')
// (8, 6, 'neigh_op_tnl_7')
// (8, 6, 'sp4_v_b_26')
// (8, 7, 'neigh_op_lft_7')
// (8, 7, 'sp4_v_b_15')
// (8, 8, 'neigh_op_bnl_7')
// (8, 8, 'sp4_v_b_2')

wire n354;
// (6, 7, 'neigh_op_tnr_0')
// (6, 8, 'neigh_op_rgt_0')
// (6, 9, 'neigh_op_bnr_0')
// (7, 7, 'neigh_op_top_0')
// (7, 8, 'lutff_0/out')
// (7, 9, 'local_g1_0')
// (7, 9, 'lutff_0/in_1')
// (7, 9, 'lutff_6/in_1')
// (7, 9, 'neigh_op_bot_0')
// (8, 7, 'neigh_op_tnl_0')
// (8, 8, 'neigh_op_lft_0')
// (8, 9, 'neigh_op_bnl_0')

wire n355;
// (6, 7, 'neigh_op_tnr_1')
// (6, 8, 'neigh_op_rgt_1')
// (6, 9, 'neigh_op_bnr_1')
// (7, 7, 'neigh_op_top_1')
// (7, 8, 'local_g1_1')
// (7, 8, 'local_g2_1')
// (7, 8, 'lutff_1/out')
// (7, 8, 'lutff_2/in_3')
// (7, 8, 'lutff_3/in_3')
// (7, 9, 'neigh_op_bot_1')
// (8, 7, 'neigh_op_tnl_1')
// (8, 8, 'local_g1_1')
// (8, 8, 'lutff_7/in_3')
// (8, 8, 'neigh_op_lft_1')
// (8, 9, 'neigh_op_bnl_1')

reg n356 = 0;
// (6, 7, 'neigh_op_tnr_2')
// (6, 8, 'local_g3_2')
// (6, 8, 'lutff_3/in_0')
// (6, 8, 'neigh_op_rgt_2')
// (6, 9, 'neigh_op_bnr_2')
// (7, 7, 'neigh_op_top_2')
// (7, 8, 'local_g0_2')
// (7, 8, 'lutff_0/in_2')
// (7, 8, 'lutff_2/out')
// (7, 9, 'neigh_op_bot_2')
// (8, 7, 'neigh_op_tnl_2')
// (8, 8, 'neigh_op_lft_2')
// (8, 9, 'neigh_op_bnl_2')

reg n357 = 0;
// (6, 7, 'neigh_op_tnr_3')
// (6, 8, 'neigh_op_rgt_3')
// (6, 9, 'neigh_op_bnr_3')
// (7, 7, 'neigh_op_top_3')
// (7, 8, 'local_g2_3')
// (7, 8, 'local_g3_3')
// (7, 8, 'lutff_2/in_1')
// (7, 8, 'lutff_3/out')
// (7, 8, 'lutff_6/in_2')
// (7, 9, 'neigh_op_bot_3')
// (8, 7, 'neigh_op_tnl_3')
// (8, 8, 'neigh_op_lft_3')
// (8, 9, 'neigh_op_bnl_3')

reg n358 = 0;
// (6, 7, 'neigh_op_tnr_4')
// (6, 8, 'neigh_op_rgt_4')
// (6, 9, 'neigh_op_bnr_4')
// (7, 7, 'neigh_op_top_4')
// (7, 8, 'local_g0_4')
// (7, 8, 'local_g1_4')
// (7, 8, 'lutff_3/in_1')
// (7, 8, 'lutff_4/out')
// (7, 8, 'lutff_7/in_2')
// (7, 9, 'neigh_op_bot_4')
// (8, 7, 'neigh_op_tnl_4')
// (8, 8, 'neigh_op_lft_4')
// (8, 9, 'neigh_op_bnl_4')

reg n359 = 0;
// (6, 7, 'neigh_op_tnr_6')
// (6, 8, 'neigh_op_rgt_6')
// (6, 9, 'neigh_op_bnr_6')
// (7, 7, 'neigh_op_top_6')
// (7, 8, 'local_g1_6')
// (7, 8, 'lutff_0/in_1')
// (7, 8, 'lutff_6/out')
// (7, 9, 'neigh_op_bot_6')
// (8, 7, 'neigh_op_tnl_6')
// (8, 8, 'neigh_op_lft_6')
// (8, 9, 'neigh_op_bnl_6')

reg n360 = 0;
// (6, 7, 'neigh_op_tnr_7')
// (6, 8, 'neigh_op_rgt_7')
// (6, 9, 'neigh_op_bnr_7')
// (7, 7, 'neigh_op_top_7')
// (7, 8, 'local_g2_7')
// (7, 8, 'lutff_6/in_1')
// (7, 8, 'lutff_7/out')
// (7, 9, 'neigh_op_bot_7')
// (8, 7, 'neigh_op_tnl_7')
// (8, 8, 'neigh_op_lft_7')
// (8, 9, 'neigh_op_bnl_7')

wire n361;
// (6, 8, 'neigh_op_tnr_0')
// (6, 9, 'neigh_op_rgt_0')
// (6, 10, 'neigh_op_bnr_0')
// (7, 8, 'neigh_op_top_0')
// (7, 9, 'local_g3_0')
// (7, 9, 'lutff_0/out')
// (7, 9, 'lutff_3/in_0')
// (7, 10, 'neigh_op_bot_0')
// (8, 8, 'neigh_op_tnl_0')
// (8, 9, 'neigh_op_lft_0')
// (8, 10, 'neigh_op_bnl_0')

wire n362;
// (6, 8, 'neigh_op_tnr_2')
// (6, 9, 'neigh_op_rgt_2')
// (6, 10, 'neigh_op_bnr_2')
// (7, 8, 'neigh_op_top_2')
// (7, 9, 'local_g0_2')
// (7, 9, 'lutff_2/out')
// (7, 9, 'lutff_3/in_1')
// (7, 10, 'neigh_op_bot_2')
// (8, 8, 'neigh_op_tnl_2')
// (8, 9, 'neigh_op_lft_2')
// (8, 10, 'neigh_op_bnl_2')

reg n363 = 0;
// (6, 8, 'neigh_op_tnr_4')
// (6, 9, 'neigh_op_rgt_4')
// (6, 10, 'neigh_op_bnr_4')
// (7, 8, 'neigh_op_top_4')
// (7, 9, 'local_g1_4')
// (7, 9, 'lutff_4/out')
// (7, 9, 'lutff_5/in_0')
// (7, 10, 'neigh_op_bot_4')
// (8, 8, 'neigh_op_tnl_4')
// (8, 9, 'neigh_op_lft_4')
// (8, 10, 'neigh_op_bnl_4')

reg n364 = 0;
// (6, 8, 'neigh_op_tnr_5')
// (6, 8, 'sp4_r_v_b_39')
// (6, 9, 'neigh_op_rgt_5')
// (6, 9, 'sp4_r_v_b_26')
// (6, 10, 'neigh_op_bnr_5')
// (6, 10, 'sp4_r_v_b_15')
// (6, 11, 'sp4_r_v_b_2')
// (7, 7, 'sp4_v_t_39')
// (7, 8, 'neigh_op_top_5')
// (7, 8, 'sp4_v_b_39')
// (7, 9, 'lutff_5/out')
// (7, 9, 'sp4_v_b_26')
// (7, 10, 'neigh_op_bot_5')
// (7, 10, 'sp4_v_b_15')
// (7, 11, 'local_g0_2')
// (7, 11, 'lutff_4/in_0')
// (7, 11, 'sp4_v_b_2')
// (8, 8, 'neigh_op_tnl_5')
// (8, 9, 'neigh_op_lft_5')
// (8, 10, 'neigh_op_bnl_5')

reg n365 = 0;
// (6, 8, 'neigh_op_tnr_6')
// (6, 9, 'neigh_op_rgt_6')
// (6, 10, 'neigh_op_bnr_6')
// (7, 8, 'neigh_op_top_6')
// (7, 9, 'local_g0_6')
// (7, 9, 'lutff_4/in_0')
// (7, 9, 'lutff_6/out')
// (7, 10, 'neigh_op_bot_6')
// (8, 8, 'neigh_op_tnl_6')
// (8, 9, 'neigh_op_lft_6')
// (8, 10, 'neigh_op_bnl_6')

reg n366 = 0;
// (6, 8, 'neigh_op_tnr_7')
// (6, 9, 'neigh_op_rgt_7')
// (6, 9, 'sp4_h_r_3')
// (6, 10, 'neigh_op_bnr_7')
// (7, 8, 'neigh_op_top_7')
// (7, 9, 'lutff_7/out')
// (7, 9, 'sp4_h_r_14')
// (7, 10, 'neigh_op_bot_7')
// (8, 8, 'neigh_op_tnl_7')
// (8, 9, 'neigh_op_lft_7')
// (8, 9, 'sp4_h_r_27')
// (8, 10, 'neigh_op_bnl_7')
// (9, 9, 'local_g2_6')
// (9, 9, 'lutff_6/in_0')
// (9, 9, 'sp4_h_r_38')
// (10, 9, 'sp4_h_l_38')

wire n367;
// (6, 9, 'neigh_op_tnr_0')
// (6, 10, 'neigh_op_rgt_0')
// (6, 11, 'neigh_op_bnr_0')
// (7, 6, 'sp12_v_t_23')
// (7, 7, 'sp12_v_b_23')
// (7, 8, 'sp12_v_b_20')
// (7, 9, 'neigh_op_top_0')
// (7, 9, 'sp12_v_b_19')
// (7, 10, 'lutff_0/out')
// (7, 10, 'sp12_v_b_16')
// (7, 11, 'neigh_op_bot_0')
// (7, 11, 'sp12_v_b_15')
// (7, 12, 'sp12_v_b_12')
// (7, 13, 'local_g3_3')
// (7, 13, 'lutff_1/in_1')
// (7, 13, 'lutff_7/in_1')
// (7, 13, 'sp12_v_b_11')
// (7, 14, 'sp12_v_b_8')
// (7, 15, 'sp12_v_b_7')
// (7, 16, 'sp12_v_b_4')
// (7, 17, 'span12_vert_3')
// (8, 9, 'neigh_op_tnl_0')
// (8, 10, 'neigh_op_lft_0')
// (8, 11, 'neigh_op_bnl_0')

wire n368;
// (6, 9, 'neigh_op_tnr_1')
// (6, 10, 'local_g2_1')
// (6, 10, 'lutff_6/in_3')
// (6, 10, 'neigh_op_rgt_1')
// (6, 11, 'neigh_op_bnr_1')
// (7, 9, 'neigh_op_top_1')
// (7, 10, 'local_g1_1')
// (7, 10, 'local_g2_1')
// (7, 10, 'lutff_1/out')
// (7, 10, 'lutff_5/in_3')
// (7, 10, 'lutff_6/in_3')
// (7, 11, 'neigh_op_bot_1')
// (8, 9, 'neigh_op_tnl_1')
// (8, 10, 'neigh_op_lft_1')
// (8, 11, 'neigh_op_bnl_1')

reg n369 = 0;
// (6, 9, 'neigh_op_tnr_2')
// (6, 10, 'neigh_op_rgt_2')
// (6, 11, 'neigh_op_bnr_2')
// (7, 9, 'neigh_op_top_2')
// (7, 10, 'local_g2_2')
// (7, 10, 'lutff_0/in_2')
// (7, 10, 'lutff_2/out')
// (7, 10, 'lutff_5/in_1')
// (7, 11, 'neigh_op_bot_2')
// (8, 9, 'neigh_op_tnl_2')
// (8, 10, 'neigh_op_lft_2')
// (8, 11, 'neigh_op_bnl_2')

reg n370 = 0;
// (6, 9, 'neigh_op_tnr_3')
// (6, 10, 'neigh_op_rgt_3')
// (6, 11, 'neigh_op_bnr_3')
// (7, 9, 'neigh_op_top_3')
// (7, 10, 'local_g0_3')
// (7, 10, 'local_g1_3')
// (7, 10, 'lutff_2/in_1')
// (7, 10, 'lutff_3/out')
// (7, 10, 'lutff_4/in_2')
// (7, 11, 'neigh_op_bot_3')
// (8, 9, 'neigh_op_tnl_3')
// (8, 10, 'neigh_op_lft_3')
// (8, 11, 'neigh_op_bnl_3')

reg n371 = 0;
// (6, 9, 'neigh_op_tnr_4')
// (6, 10, 'neigh_op_rgt_4')
// (6, 11, 'neigh_op_bnr_4')
// (7, 9, 'neigh_op_top_4')
// (7, 10, 'local_g1_4')
// (7, 10, 'lutff_0/in_1')
// (7, 10, 'lutff_4/out')
// (7, 11, 'neigh_op_bot_4')
// (8, 9, 'neigh_op_tnl_4')
// (8, 10, 'neigh_op_lft_4')
// (8, 11, 'neigh_op_bnl_4')

reg n372 = 0;
// (6, 9, 'neigh_op_tnr_6')
// (6, 10, 'neigh_op_rgt_6')
// (6, 11, 'neigh_op_bnr_6')
// (7, 9, 'neigh_op_top_6')
// (7, 10, 'local_g2_6')
// (7, 10, 'local_g3_6')
// (7, 10, 'lutff_3/in_1')
// (7, 10, 'lutff_6/out')
// (7, 10, 'lutff_7/in_2')
// (7, 11, 'neigh_op_bot_6')
// (8, 9, 'neigh_op_tnl_6')
// (8, 10, 'neigh_op_lft_6')
// (8, 11, 'neigh_op_bnl_6')

reg n373 = 0;
// (6, 9, 'neigh_op_tnr_7')
// (6, 10, 'neigh_op_rgt_7')
// (6, 11, 'neigh_op_bnr_7')
// (7, 9, 'neigh_op_top_7')
// (7, 10, 'local_g0_7')
// (7, 10, 'lutff_4/in_1')
// (7, 10, 'lutff_7/out')
// (7, 11, 'neigh_op_bot_7')
// (8, 9, 'neigh_op_tnl_7')
// (8, 10, 'neigh_op_lft_7')
// (8, 11, 'neigh_op_bnl_7')

reg n374 = 0;
// (6, 9, 'sp12_h_r_0')
// (7, 9, 'sp12_h_r_3')
// (8, 9, 'sp12_h_r_4')
// (9, 9, 'local_g0_7')
// (9, 9, 'lutff_3/in_0')
// (9, 9, 'sp12_h_r_7')
// (10, 9, 'sp12_h_r_8')
// (11, 8, 'neigh_op_tnr_2')
// (11, 9, 'neigh_op_rgt_2')
// (11, 9, 'sp12_h_r_11')
// (11, 10, 'neigh_op_bnr_2')
// (12, 8, 'neigh_op_top_2')
// (12, 9, 'lutff_2/out')
// (12, 9, 'sp12_h_r_12')
// (12, 10, 'neigh_op_bot_2')
// (13, 8, 'logic_op_tnl_2')
// (13, 9, 'logic_op_lft_2')
// (13, 9, 'span12_horz_12')
// (13, 10, 'logic_op_bnl_2')

wire \d_out[4] ;
// (6, 9, 'sp12_h_r_1')
// (7, 9, 'sp12_h_r_2')
// (8, 9, 'sp12_h_r_5')
// (9, 9, 'sp12_h_r_6')
// (10, 8, 'neigh_op_tnr_1')
// (10, 9, 'neigh_op_rgt_1')
// (10, 9, 'sp12_h_r_9')
// (10, 10, 'neigh_op_bnr_1')
// (11, 8, 'neigh_op_top_1')
// (11, 9, 'lutff_1/out')
// (11, 9, 'sp12_h_r_10')
// (11, 10, 'neigh_op_bot_1')
// (12, 8, 'neigh_op_tnl_1')
// (12, 9, 'neigh_op_lft_1')
// (12, 9, 'sp12_h_r_13')
// (12, 10, 'neigh_op_bnl_1')
// (13, 9, 'io_1/D_OUT_0')
// (13, 9, 'io_1/PAD')
// (13, 9, 'local_g0_5')
// (13, 9, 'span12_horz_13')

wire n376;
// (6, 10, 'neigh_op_tnr_0')
// (6, 11, 'neigh_op_rgt_0')
// (6, 12, 'neigh_op_bnr_0')
// (7, 0, 'span12_vert_20')
// (7, 1, 'sp12_v_b_20')
// (7, 2, 'sp12_v_b_19')
// (7, 3, 'sp12_v_b_16')
// (7, 4, 'sp12_v_b_15')
// (7, 5, 'sp12_v_b_12')
// (7, 6, 'sp12_v_b_11')
// (7, 7, 'sp12_v_b_8')
// (7, 8, 'sp12_v_b_7')
// (7, 9, 'local_g3_4')
// (7, 9, 'lutff_2/in_3')
// (7, 9, 'sp12_v_b_4')
// (7, 10, 'neigh_op_top_0')
// (7, 10, 'sp12_v_b_3')
// (7, 11, 'lutff_0/out')
// (7, 11, 'sp12_v_b_0')
// (7, 12, 'neigh_op_bot_0')
// (8, 10, 'neigh_op_tnl_0')
// (8, 11, 'neigh_op_lft_0')
// (8, 12, 'neigh_op_bnl_0')

reg n377 = 0;
// (6, 10, 'neigh_op_tnr_1')
// (6, 11, 'neigh_op_rgt_1')
// (6, 12, 'neigh_op_bnr_1')
// (7, 10, 'neigh_op_top_1')
// (7, 11, 'local_g0_1')
// (7, 11, 'lutff_1/out')
// (7, 11, 'lutff_3/in_0')
// (7, 12, 'neigh_op_bot_1')
// (8, 10, 'neigh_op_tnl_1')
// (8, 11, 'neigh_op_lft_1')
// (8, 12, 'neigh_op_bnl_1')

reg n378 = 0;
// (6, 10, 'neigh_op_tnr_3')
// (6, 11, 'neigh_op_rgt_3')
// (6, 12, 'neigh_op_bnr_3')
// (7, 10, 'neigh_op_top_3')
// (7, 11, 'local_g1_3')
// (7, 11, 'lutff_2/in_0')
// (7, 11, 'lutff_3/out')
// (7, 12, 'neigh_op_bot_3')
// (8, 10, 'neigh_op_tnl_3')
// (8, 11, 'neigh_op_lft_3')
// (8, 12, 'neigh_op_bnl_3')

reg n379 = 0;
// (6, 10, 'neigh_op_tnr_4')
// (6, 11, 'neigh_op_rgt_4')
// (6, 12, 'neigh_op_bnr_4')
// (7, 10, 'neigh_op_top_4')
// (7, 11, 'local_g0_4')
// (7, 11, 'local_g1_4')
// (7, 11, 'lutff_0/in_1')
// (7, 11, 'lutff_4/out')
// (7, 11, 'lutff_7/in_1')
// (7, 12, 'neigh_op_bot_4')
// (8, 10, 'neigh_op_tnl_4')
// (8, 11, 'neigh_op_lft_4')
// (8, 12, 'neigh_op_bnl_4')

reg n380 = 0;
// (6, 10, 'neigh_op_tnr_6')
// (6, 11, 'neigh_op_rgt_6')
// (6, 12, 'neigh_op_bnr_6')
// (7, 10, 'neigh_op_top_6')
// (7, 11, 'lutff_6/out')
// (7, 12, 'neigh_op_bot_6')
// (8, 10, 'local_g3_6')
// (8, 10, 'lutff_3/in_0')
// (8, 10, 'neigh_op_tnl_6')
// (8, 11, 'neigh_op_lft_6')
// (8, 12, 'neigh_op_bnl_6')

reg n381 = 0;
// (6, 10, 'neigh_op_tnr_7')
// (6, 11, 'neigh_op_rgt_7')
// (6, 12, 'neigh_op_bnr_7')
// (7, 10, 'neigh_op_top_7')
// (7, 11, 'local_g2_7')
// (7, 11, 'lutff_1/in_0')
// (7, 11, 'lutff_7/out')
// (7, 12, 'neigh_op_bot_7')
// (8, 10, 'neigh_op_tnl_7')
// (8, 11, 'neigh_op_lft_7')
// (8, 12, 'neigh_op_bnl_7')

reg n382 = 0;
// (6, 11, 'neigh_op_tnr_3')
// (6, 12, 'neigh_op_rgt_3')
// (6, 13, 'neigh_op_bnr_3')
// (7, 11, 'neigh_op_top_3')
// (7, 12, 'local_g1_3')
// (7, 12, 'lutff_3/out')
// (7, 12, 'lutff_4/in_0')
// (7, 13, 'neigh_op_bot_3')
// (8, 11, 'neigh_op_tnl_3')
// (8, 12, 'neigh_op_lft_3')
// (8, 13, 'neigh_op_bnl_3')

reg n383 = 0;
// (6, 11, 'neigh_op_tnr_4')
// (6, 12, 'neigh_op_rgt_4')
// (6, 13, 'neigh_op_bnr_4')
// (7, 11, 'neigh_op_top_4')
// (7, 12, 'local_g1_4')
// (7, 12, 'lutff_1/in_0')
// (7, 12, 'lutff_4/out')
// (7, 13, 'neigh_op_bot_4')
// (8, 11, 'neigh_op_tnl_4')
// (8, 12, 'neigh_op_lft_4')
// (8, 13, 'neigh_op_bnl_4')

reg n384 = 0;
// (6, 11, 'neigh_op_tnr_5')
// (6, 12, 'neigh_op_rgt_5')
// (6, 13, 'neigh_op_bnr_5')
// (7, 11, 'neigh_op_top_5')
// (7, 12, 'local_g0_5')
// (7, 12, 'lutff_5/out')
// (7, 12, 'lutff_7/in_0')
// (7, 13, 'neigh_op_bot_5')
// (8, 11, 'neigh_op_tnl_5')
// (8, 12, 'neigh_op_lft_5')
// (8, 13, 'neigh_op_bnl_5')

reg n385 = 0;
// (6, 11, 'neigh_op_tnr_6')
// (6, 11, 'sp4_r_v_b_41')
// (6, 12, 'neigh_op_rgt_6')
// (6, 12, 'sp4_r_v_b_28')
// (6, 13, 'neigh_op_bnr_6')
// (6, 13, 'sp4_r_v_b_17')
// (6, 14, 'sp4_r_v_b_4')
// (7, 10, 'sp4_v_t_41')
// (7, 11, 'neigh_op_top_6')
// (7, 11, 'sp4_v_b_41')
// (7, 12, 'lutff_6/out')
// (7, 12, 'sp4_v_b_28')
// (7, 13, 'neigh_op_bot_6')
// (7, 13, 'sp4_v_b_17')
// (7, 14, 'local_g1_4')
// (7, 14, 'lutff_7/in_0')
// (7, 14, 'sp4_v_b_4')
// (8, 11, 'neigh_op_tnl_6')
// (8, 12, 'neigh_op_lft_6')
// (8, 13, 'neigh_op_bnl_6')

reg n386 = 0;
// (6, 11, 'neigh_op_tnr_7')
// (6, 12, 'neigh_op_rgt_7')
// (6, 13, 'neigh_op_bnr_7')
// (7, 11, 'neigh_op_top_7')
// (7, 12, 'local_g1_7')
// (7, 12, 'lutff_6/in_0')
// (7, 12, 'lutff_7/out')
// (7, 13, 'neigh_op_bot_7')
// (8, 11, 'neigh_op_tnl_7')
// (8, 12, 'neigh_op_lft_7')
// (8, 13, 'neigh_op_bnl_7')

wire n387;
// (6, 11, 'sp4_r_v_b_37')
// (6, 12, 'sp4_r_v_b_24')
// (6, 13, 'neigh_op_tnr_0')
// (6, 13, 'sp4_r_v_b_13')
// (6, 14, 'neigh_op_rgt_0')
// (6, 14, 'sp4_r_v_b_0')
// (6, 15, 'neigh_op_bnr_0')
// (7, 10, 'sp4_v_t_37')
// (7, 11, 'sp4_v_b_37')
// (7, 12, 'sp4_v_b_24')
// (7, 13, 'local_g0_5')
// (7, 13, 'lutff_0/in_3')
// (7, 13, 'neigh_op_top_0')
// (7, 13, 'sp4_v_b_13')
// (7, 14, 'lutff_0/out')
// (7, 14, 'sp4_v_b_0')
// (7, 15, 'neigh_op_bot_0')
// (8, 13, 'neigh_op_tnl_0')
// (8, 14, 'neigh_op_lft_0')
// (8, 15, 'neigh_op_bnl_0')

wire n388;
// (6, 12, 'neigh_op_tnr_0')
// (6, 13, 'neigh_op_rgt_0')
// (6, 14, 'neigh_op_bnr_0')
// (7, 12, 'local_g1_0')
// (7, 12, 'lutff_0/in_3')
// (7, 12, 'neigh_op_top_0')
// (7, 13, 'lutff_0/out')
// (7, 14, 'neigh_op_bot_0')
// (8, 12, 'neigh_op_tnl_0')
// (8, 13, 'neigh_op_lft_0')
// (8, 14, 'neigh_op_bnl_0')

wire n389;
// (6, 12, 'neigh_op_tnr_4')
// (6, 13, 'neigh_op_rgt_4')
// (6, 14, 'neigh_op_bnr_4')
// (7, 12, 'neigh_op_top_4')
// (7, 13, 'local_g0_4')
// (7, 13, 'lutff_4/out')
// (7, 13, 'lutff_5/in_3')
// (7, 14, 'neigh_op_bot_4')
// (8, 12, 'neigh_op_tnl_4')
// (8, 13, 'neigh_op_lft_4')
// (8, 14, 'neigh_op_bnl_4')

wire n390;
// (6, 12, 'neigh_op_tnr_5')
// (6, 13, 'neigh_op_rgt_5')
// (6, 14, 'neigh_op_bnr_5')
// (7, 12, 'neigh_op_top_5')
// (7, 13, 'local_g1_5')
// (7, 13, 'lutff_1/in_3')
// (7, 13, 'lutff_5/out')
// (7, 14, 'neigh_op_bot_5')
// (8, 12, 'neigh_op_tnl_5')
// (8, 13, 'neigh_op_lft_5')
// (8, 14, 'neigh_op_bnl_5')

reg n391 = 0;
// (6, 12, 'neigh_op_tnr_7')
// (6, 13, 'neigh_op_rgt_7')
// (6, 14, 'neigh_op_bnr_7')
// (7, 12, 'neigh_op_top_7')
// (7, 13, 'lutff_7/out')
// (7, 14, 'neigh_op_bot_7')
// (8, 12, 'neigh_op_tnl_7')
// (8, 13, 'local_g0_7')
// (8, 13, 'lutff_7/in_0')
// (8, 13, 'neigh_op_lft_7')
// (8, 14, 'neigh_op_bnl_7')

reg n392 = 0;
// (6, 12, 'sp4_h_r_11')
// (7, 12, 'local_g0_6')
// (7, 12, 'local_g1_6')
// (7, 12, 'lutff_0/in_2')
// (7, 12, 'lutff_5/in_2')
// (7, 12, 'sp4_h_r_22')
// (8, 6, 'neigh_op_tnr_3')
// (8, 7, 'neigh_op_rgt_3')
// (8, 8, 'neigh_op_bnr_3')
// (8, 12, 'sp4_h_r_35')
// (9, 4, 'sp4_r_v_b_42')
// (9, 5, 'local_g0_7')
// (9, 5, 'lutff_7/in_0')
// (9, 5, 'sp4_r_v_b_31')
// (9, 5, 'sp4_r_v_b_47')
// (9, 6, 'neigh_op_top_3')
// (9, 6, 'sp12_v_t_22')
// (9, 6, 'sp4_r_v_b_18')
// (9, 6, 'sp4_r_v_b_34')
// (9, 7, 'lutff_3/out')
// (9, 7, 'sp12_v_b_22')
// (9, 7, 'sp4_r_v_b_23')
// (9, 7, 'sp4_r_v_b_7')
// (9, 8, 'neigh_op_bot_3')
// (9, 8, 'sp12_v_b_21')
// (9, 8, 'sp4_r_v_b_10')
// (9, 9, 'sp12_v_b_18')
// (9, 9, 'sp4_r_v_b_43')
// (9, 10, 'sp12_v_b_17')
// (9, 10, 'sp4_r_v_b_30')
// (9, 11, 'sp12_v_b_14')
// (9, 11, 'sp4_r_v_b_19')
// (9, 12, 'local_g2_5')
// (9, 12, 'lutff_5/in_0')
// (9, 12, 'sp12_v_b_13')
// (9, 12, 'sp4_h_r_46')
// (9, 12, 'sp4_r_v_b_6')
// (9, 13, 'sp12_v_b_10')
// (9, 14, 'sp12_v_b_9')
// (9, 15, 'sp12_v_b_6')
// (9, 16, 'sp12_v_b_5')
// (9, 17, 'span12_vert_2')
// (10, 3, 'sp4_v_t_42')
// (10, 4, 'sp4_v_b_42')
// (10, 4, 'sp4_v_t_47')
// (10, 5, 'sp4_v_b_31')
// (10, 5, 'sp4_v_b_47')
// (10, 6, 'neigh_op_tnl_3')
// (10, 6, 'sp4_v_b_18')
// (10, 6, 'sp4_v_b_34')
// (10, 7, 'neigh_op_lft_3')
// (10, 7, 'sp4_v_b_23')
// (10, 7, 'sp4_v_b_7')
// (10, 8, 'neigh_op_bnl_3')
// (10, 8, 'sp4_v_b_10')
// (10, 8, 'sp4_v_t_43')
// (10, 9, 'sp4_v_b_43')
// (10, 10, 'sp4_v_b_30')
// (10, 11, 'sp4_v_b_19')
// (10, 12, 'sp4_h_l_46')
// (10, 12, 'sp4_v_b_6')

reg n393 = 0;
// (6, 13, 'neigh_op_tnr_3')
// (6, 14, 'neigh_op_rgt_3')
// (6, 15, 'neigh_op_bnr_3')
// (7, 13, 'neigh_op_top_3')
// (7, 14, 'local_g0_3')
// (7, 14, 'lutff_3/out')
// (7, 14, 'lutff_5/in_0')
// (7, 15, 'neigh_op_bot_3')
// (8, 13, 'neigh_op_tnl_3')
// (8, 14, 'neigh_op_lft_3')
// (8, 15, 'neigh_op_bnl_3')

reg n394 = 0;
// (6, 13, 'neigh_op_tnr_5')
// (6, 14, 'neigh_op_rgt_5')
// (6, 15, 'neigh_op_bnr_5')
// (7, 13, 'neigh_op_top_5')
// (7, 14, 'lutff_5/out')
// (7, 14, 'sp4_r_v_b_43')
// (7, 15, 'local_g0_6')
// (7, 15, 'lutff_2/in_0')
// (7, 15, 'neigh_op_bot_5')
// (7, 15, 'sp4_r_v_b_30')
// (7, 16, 'sp4_r_v_b_19')
// (8, 13, 'neigh_op_tnl_5')
// (8, 13, 'sp4_v_t_43')
// (8, 14, 'neigh_op_lft_5')
// (8, 14, 'sp4_v_b_43')
// (8, 15, 'neigh_op_bnl_5')
// (8, 15, 'sp4_v_b_30')
// (8, 16, 'sp4_v_b_19')
// (8, 17, 'span4_vert_6')

reg n395 = 0;
// (6, 13, 'neigh_op_tnr_7')
// (6, 14, 'neigh_op_rgt_7')
// (6, 15, 'neigh_op_bnr_7')
// (7, 13, 'neigh_op_top_7')
// (7, 14, 'local_g0_7')
// (7, 14, 'local_g1_7')
// (7, 14, 'lutff_0/in_1')
// (7, 14, 'lutff_3/in_1')
// (7, 14, 'lutff_7/out')
// (7, 15, 'neigh_op_bot_7')
// (8, 13, 'neigh_op_tnl_7')
// (8, 14, 'neigh_op_lft_7')
// (8, 15, 'neigh_op_bnl_7')

reg n396 = 0;
// (6, 14, 'neigh_op_tnr_0')
// (6, 15, 'neigh_op_rgt_0')
// (6, 16, 'neigh_op_bnr_0')
// (7, 14, 'neigh_op_top_0')
// (7, 15, 'local_g1_0')
// (7, 15, 'lutff_0/out')
// (7, 15, 'lutff_1/in_0')
// (7, 16, 'neigh_op_bot_0')
// (8, 14, 'neigh_op_tnl_0')
// (8, 15, 'neigh_op_lft_0')
// (8, 16, 'neigh_op_bnl_0')

reg n397 = 0;
// (6, 14, 'neigh_op_tnr_1')
// (6, 15, 'neigh_op_rgt_1')
// (6, 16, 'neigh_op_bnr_1')
// (7, 4, 'sp12_v_t_22')
// (7, 5, 'sp12_v_b_22')
// (7, 6, 'sp12_v_b_21')
// (7, 7, 'sp12_v_b_18')
// (7, 8, 'sp12_v_b_17')
// (7, 9, 'sp12_v_b_14')
// (7, 10, 'sp12_v_b_13')
// (7, 11, 'sp12_v_b_10')
// (7, 12, 'local_g2_1')
// (7, 12, 'lutff_5/in_0')
// (7, 12, 'sp12_v_b_9')
// (7, 13, 'local_g2_6')
// (7, 13, 'lutff_0/in_0')
// (7, 13, 'sp12_v_b_6')
// (7, 14, 'local_g0_1')
// (7, 14, 'lutff_3/in_0')
// (7, 14, 'neigh_op_top_1')
// (7, 14, 'sp12_v_b_5')
// (7, 15, 'local_g0_1')
// (7, 15, 'lutff_1/out')
// (7, 15, 'lutff_3/in_0')
// (7, 15, 'sp12_v_b_2')
// (7, 16, 'neigh_op_bot_1')
// (7, 16, 'sp12_v_b_1')
// (8, 14, 'neigh_op_tnl_1')
// (8, 15, 'neigh_op_lft_1')
// (8, 16, 'neigh_op_bnl_1')

reg n398 = 0;
// (6, 14, 'neigh_op_tnr_2')
// (6, 15, 'neigh_op_rgt_2')
// (6, 16, 'neigh_op_bnr_2')
// (7, 14, 'neigh_op_top_2')
// (7, 15, 'local_g1_2')
// (7, 15, 'lutff_2/out')
// (7, 15, 'lutff_5/in_0')
// (7, 16, 'neigh_op_bot_2')
// (8, 14, 'neigh_op_tnl_2')
// (8, 15, 'neigh_op_lft_2')
// (8, 16, 'neigh_op_bnl_2')

reg n399 = 0;
// (6, 14, 'neigh_op_tnr_3')
// (6, 15, 'neigh_op_rgt_3')
// (6, 16, 'neigh_op_bnr_3')
// (7, 14, 'neigh_op_top_3')
// (7, 15, 'local_g0_3')
// (7, 15, 'lutff_3/out')
// (7, 15, 'lutff_7/in_0')
// (7, 16, 'neigh_op_bot_3')
// (8, 14, 'neigh_op_tnl_3')
// (8, 15, 'neigh_op_lft_3')
// (8, 16, 'neigh_op_bnl_3')

reg n400 = 0;
// (6, 14, 'neigh_op_tnr_5')
// (6, 15, 'neigh_op_rgt_5')
// (6, 16, 'neigh_op_bnr_5')
// (7, 14, 'local_g1_5')
// (7, 14, 'lutff_0/in_0')
// (7, 14, 'neigh_op_top_5')
// (7, 15, 'local_g1_5')
// (7, 15, 'lutff_3/in_1')
// (7, 15, 'lutff_5/out')
// (7, 16, 'neigh_op_bot_5')
// (8, 14, 'neigh_op_tnl_5')
// (8, 15, 'neigh_op_lft_5')
// (8, 16, 'neigh_op_bnl_5')

reg n401 = 0;
// (6, 14, 'neigh_op_tnr_7')
// (6, 15, 'neigh_op_rgt_7')
// (6, 16, 'neigh_op_bnr_7')
// (7, 14, 'neigh_op_top_7')
// (7, 15, 'local_g1_7')
// (7, 15, 'lutff_0/in_0')
// (7, 15, 'lutff_7/out')
// (7, 16, 'neigh_op_bot_7')
// (8, 14, 'neigh_op_tnl_7')
// (8, 15, 'neigh_op_lft_7')
// (8, 16, 'neigh_op_bnl_7')

wire n402;
// (7, 1, 'neigh_op_tnr_0')
// (7, 1, 'sp4_r_v_b_29')
// (7, 2, 'local_g2_0')
// (7, 2, 'local_g3_0')
// (7, 2, 'lutff_1/in_2')
// (7, 2, 'lutff_7/in_1')
// (7, 2, 'neigh_op_rgt_0')
// (7, 2, 'sp4_r_v_b_16')
// (7, 3, 'local_g1_0')
// (7, 3, 'local_g1_5')
// (7, 3, 'lutff_0/in_3')
// (7, 3, 'lutff_3/in_3')
// (7, 3, 'neigh_op_bnr_0')
// (7, 3, 'sp4_r_v_b_5')
// (8, 0, 'span4_vert_29')
// (8, 1, 'neigh_op_top_0')
// (8, 1, 'sp4_v_b_29')
// (8, 2, 'local_g1_0')
// (8, 2, 'lutff_0/out')
// (8, 2, 'lutff_6/in_1')
// (8, 2, 'sp4_v_b_16')
// (8, 3, 'neigh_op_bot_0')
// (8, 3, 'sp4_v_b_5')
// (9, 1, 'neigh_op_tnl_0')
// (9, 2, 'neigh_op_lft_0')
// (9, 3, 'neigh_op_bnl_0')

wire n403;
// (7, 1, 'neigh_op_tnr_3')
// (7, 2, 'local_g3_3')
// (7, 2, 'lutff_3/in_3')
// (7, 2, 'neigh_op_rgt_3')
// (7, 3, 'neigh_op_bnr_3')
// (8, 1, 'neigh_op_top_3')
// (8, 2, 'lutff_3/out')
// (8, 3, 'neigh_op_bot_3')
// (9, 1, 'neigh_op_tnl_3')
// (9, 2, 'neigh_op_lft_3')
// (9, 3, 'neigh_op_bnl_3')

wire n404;
// (7, 1, 'sp4_r_v_b_25')
// (7, 1, 'sp4_r_v_b_30')
// (7, 2, 'sp4_r_v_b_12')
// (7, 2, 'sp4_r_v_b_19')
// (7, 3, 'neigh_op_tnr_3')
// (7, 3, 'sp4_r_v_b_1')
// (7, 3, 'sp4_r_v_b_6')
// (7, 4, 'local_g2_3')
// (7, 4, 'local_g2_6')
// (7, 4, 'lutff_0/in_1')
// (7, 4, 'lutff_5/in_3')
// (7, 4, 'neigh_op_rgt_3')
// (7, 4, 'sp4_r_v_b_38')
// (7, 5, 'neigh_op_bnr_3')
// (7, 5, 'sp4_r_v_b_27')
// (7, 6, 'sp4_r_v_b_14')
// (7, 7, 'sp4_r_v_b_3')
// (8, 0, 'span4_vert_25')
// (8, 0, 'span4_vert_30')
// (8, 1, 'sp4_v_b_25')
// (8, 1, 'sp4_v_b_30')
// (8, 2, 'local_g0_3')
// (8, 2, 'lutff_0/in_1')
// (8, 2, 'sp4_v_b_12')
// (8, 2, 'sp4_v_b_19')
// (8, 3, 'local_g1_1')
// (8, 3, 'lutff_1/in_3')
// (8, 3, 'lutff_2/in_2')
// (8, 3, 'neigh_op_top_3')
// (8, 3, 'sp4_h_r_8')
// (8, 3, 'sp4_v_b_1')
// (8, 3, 'sp4_v_b_6')
// (8, 3, 'sp4_v_t_38')
// (8, 4, 'lutff_3/out')
// (8, 4, 'sp4_v_b_38')
// (8, 5, 'neigh_op_bot_3')
// (8, 5, 'sp4_v_b_27')
// (8, 6, 'sp4_v_b_14')
// (8, 7, 'sp4_v_b_3')
// (9, 3, 'neigh_op_tnl_3')
// (9, 3, 'sp4_h_r_21')
// (9, 4, 'neigh_op_lft_3')
// (9, 5, 'neigh_op_bnl_3')
// (10, 3, 'sp4_h_r_32')
// (11, 3, 'sp4_h_r_45')
// (12, 3, 'sp4_h_l_45')

wire n405;
// (7, 1, 'sp4_r_v_b_26')
// (7, 2, 'neigh_op_tnr_1')
// (7, 2, 'sp4_r_v_b_15')
// (7, 3, 'neigh_op_rgt_1')
// (7, 3, 'sp4_r_v_b_2')
// (7, 4, 'neigh_op_bnr_1')
// (8, 0, 'span4_vert_26')
// (8, 1, 'sp4_v_b_26')
// (8, 2, 'local_g0_7')
// (8, 2, 'lutff_6/in_3')
// (8, 2, 'neigh_op_top_1')
// (8, 2, 'sp4_v_b_15')
// (8, 3, 'lutff_1/out')
// (8, 3, 'sp4_v_b_2')
// (8, 4, 'neigh_op_bot_1')
// (9, 2, 'neigh_op_tnl_1')
// (9, 3, 'neigh_op_lft_1')
// (9, 4, 'neigh_op_bnl_1')

wire n406;
// (7, 1, 'sp4_r_v_b_33')
// (7, 2, 'sp4_r_v_b_20')
// (7, 3, 'sp4_r_v_b_9')
// (7, 4, 'neigh_op_tnr_5')
// (7, 5, 'neigh_op_rgt_5')
// (7, 6, 'neigh_op_bnr_5')
// (8, 0, 'span12_vert_18')
// (8, 0, 'span4_vert_33')
// (8, 1, 'sp12_v_b_18')
// (8, 1, 'sp4_v_b_33')
// (8, 2, 'sp12_v_b_17')
// (8, 2, 'sp4_r_v_b_46')
// (8, 2, 'sp4_v_b_20')
// (8, 3, 'local_g0_0')
// (8, 3, 'local_g0_1')
// (8, 3, 'lutff_5/in_1')
// (8, 3, 'lutff_7/in_2')
// (8, 3, 'sp12_v_b_14')
// (8, 3, 'sp4_r_v_b_35')
// (8, 3, 'sp4_v_b_9')
// (8, 4, 'local_g1_5')
// (8, 4, 'lutff_3/in_3')
// (8, 4, 'neigh_op_top_5')
// (8, 4, 'sp12_v_b_13')
// (8, 4, 'sp4_r_v_b_22')
// (8, 5, 'lutff_5/out')
// (8, 5, 'sp12_v_b_10')
// (8, 5, 'sp4_r_v_b_11')
// (8, 6, 'neigh_op_bot_5')
// (8, 6, 'sp12_v_b_9')
// (8, 7, 'sp12_v_b_6')
// (8, 8, 'sp12_v_b_5')
// (8, 9, 'sp12_v_b_2')
// (8, 10, 'sp12_v_b_1')
// (9, 1, 'sp4_v_t_46')
// (9, 2, 'sp4_v_b_46')
// (9, 3, 'local_g2_3')
// (9, 3, 'lutff_7/in_2')
// (9, 3, 'sp4_v_b_35')
// (9, 4, 'neigh_op_tnl_5')
// (9, 4, 'sp4_v_b_22')
// (9, 5, 'neigh_op_lft_5')
// (9, 5, 'sp4_v_b_11')
// (9, 6, 'neigh_op_bnl_5')

wire n407;
// (7, 1, 'sp4_r_v_b_34')
// (7, 2, 'local_g3_7')
// (7, 2, 'lutff_1/in_1')
// (7, 2, 'neigh_op_tnr_5')
// (7, 2, 'sp4_r_v_b_23')
// (7, 3, 'local_g3_5')
// (7, 3, 'lutff_4/in_2')
// (7, 3, 'lutff_7/in_1')
// (7, 3, 'neigh_op_rgt_5')
// (7, 3, 'sp4_r_v_b_10')
// (7, 4, 'neigh_op_bnr_5')
// (8, 0, 'span4_vert_34')
// (8, 1, 'sp4_v_b_34')
// (8, 2, 'local_g0_5')
// (8, 2, 'local_g1_5')
// (8, 2, 'lutff_0/in_2')
// (8, 2, 'lutff_1/in_3')
// (8, 2, 'lutff_3/in_3')
// (8, 2, 'lutff_5/in_2')
// (8, 2, 'neigh_op_top_5')
// (8, 2, 'sp4_v_b_23')
// (8, 3, 'lutff_5/out')
// (8, 3, 'sp4_v_b_10')
// (8, 4, 'neigh_op_bot_5')
// (9, 2, 'neigh_op_tnl_5')
// (9, 3, 'neigh_op_lft_5')
// (9, 4, 'neigh_op_bnl_5')

wire n408;
// (7, 1, 'sp4_r_v_b_39')
// (7, 2, 'local_g0_2')
// (7, 2, 'lutff_1/in_3')
// (7, 2, 'sp4_r_v_b_26')
// (7, 3, 'local_g2_1')
// (7, 3, 'local_g3_1')
// (7, 3, 'lutff_0/in_2')
// (7, 3, 'lutff_3/in_2')
// (7, 3, 'neigh_op_tnr_1')
// (7, 3, 'sp4_r_v_b_15')
// (7, 4, 'neigh_op_rgt_1')
// (7, 4, 'sp4_r_v_b_2')
// (7, 5, 'neigh_op_bnr_1')
// (8, 0, 'span4_vert_39')
// (8, 1, 'sp4_v_b_39')
// (8, 2, 'local_g3_2')
// (8, 2, 'lutff_1/in_2')
// (8, 2, 'lutff_3/in_0')
// (8, 2, 'sp4_v_b_26')
// (8, 3, 'neigh_op_top_1')
// (8, 3, 'sp4_v_b_15')
// (8, 4, 'lutff_1/out')
// (8, 4, 'sp4_v_b_2')
// (8, 5, 'neigh_op_bot_1')
// (9, 3, 'neigh_op_tnl_1')
// (9, 4, 'neigh_op_lft_1')
// (9, 5, 'neigh_op_bnl_1')

wire n409;
// (7, 1, 'sp4_r_v_b_43')
// (7, 2, 'sp4_r_v_b_30')
// (7, 3, 'sp4_r_v_b_19')
// (7, 4, 'sp4_r_v_b_6')
// (8, 0, 'span4_vert_43')
// (8, 1, 'sp4_v_b_43')
// (8, 2, 'sp4_v_b_30')
// (8, 3, 'sp4_v_b_19')
// (8, 4, 'local_g1_1')
// (8, 4, 'lutff_2/in_2')
// (8, 4, 'lutff_5/in_3')
// (8, 4, 'sp4_h_r_1')
// (8, 4, 'sp4_h_r_6')
// (8, 4, 'sp4_v_b_6')
// (9, 4, 'local_g0_3')
// (9, 4, 'lutff_0/in_3')
// (9, 4, 'sp4_h_r_12')
// (9, 4, 'sp4_h_r_19')
// (10, 3, 'neigh_op_tnr_2')
// (10, 4, 'neigh_op_rgt_2')
// (10, 4, 'sp4_h_r_25')
// (10, 4, 'sp4_h_r_30')
// (10, 5, 'neigh_op_bnr_2')
// (11, 3, 'neigh_op_top_2')
// (11, 4, 'lutff_2/out')
// (11, 4, 'sp4_h_r_36')
// (11, 4, 'sp4_h_r_43')
// (11, 5, 'neigh_op_bot_2')
// (12, 3, 'neigh_op_tnl_2')
// (12, 4, 'neigh_op_lft_2')
// (12, 4, 'sp4_h_l_36')
// (12, 4, 'sp4_h_l_43')
// (12, 5, 'neigh_op_bnl_2')

wire n410;
// (7, 2, 'local_g2_7')
// (7, 2, 'lutff_0/in_3')
// (7, 2, 'lutff_7/in_2')
// (7, 2, 'neigh_op_tnr_7')
// (7, 3, 'local_g2_7')
// (7, 3, 'lutff_2/in_1')
// (7, 3, 'neigh_op_rgt_7')
// (7, 4, 'neigh_op_bnr_7')
// (8, 2, 'neigh_op_top_7')
// (8, 3, 'lutff_7/out')
// (8, 4, 'neigh_op_bot_7')
// (9, 2, 'neigh_op_tnl_7')
// (9, 3, 'neigh_op_lft_7')
// (9, 4, 'neigh_op_bnl_7')

wire n411;
// (7, 2, 'neigh_op_tnr_0')
// (7, 3, 'local_g2_0')
// (7, 3, 'lutff_5/in_3')
// (7, 3, 'neigh_op_rgt_0')
// (7, 4, 'neigh_op_bnr_0')
// (8, 2, 'neigh_op_top_0')
// (8, 3, 'lutff_0/out')
// (8, 4, 'neigh_op_bot_0')
// (9, 2, 'neigh_op_tnl_0')
// (9, 3, 'neigh_op_lft_0')
// (9, 4, 'neigh_op_bnl_0')

wire n412;
// (7, 2, 'neigh_op_tnr_2')
// (7, 3, 'neigh_op_rgt_2')
// (7, 4, 'neigh_op_bnr_2')
// (8, 2, 'local_g0_2')
// (8, 2, 'lutff_7/in_3')
// (8, 2, 'neigh_op_top_2')
// (8, 3, 'lutff_2/out')
// (8, 4, 'neigh_op_bot_2')
// (9, 2, 'neigh_op_tnl_2')
// (9, 3, 'neigh_op_lft_2')
// (9, 4, 'neigh_op_bnl_2')

wire n413;
// (7, 2, 'neigh_op_tnr_3')
// (7, 3, 'neigh_op_rgt_3')
// (7, 4, 'neigh_op_bnr_3')
// (8, 2, 'neigh_op_top_3')
// (8, 3, 'local_g1_3')
// (8, 3, 'local_g2_3')
// (8, 3, 'lutff_0/in_3')
// (8, 3, 'lutff_1/in_0')
// (8, 3, 'lutff_2/in_0')
// (8, 3, 'lutff_3/out')
// (8, 3, 'lutff_6/in_2')
// (8, 4, 'neigh_op_bot_3')
// (9, 2, 'neigh_op_tnl_3')
// (9, 3, 'neigh_op_lft_3')
// (9, 4, 'neigh_op_bnl_3')

wire n414;
// (7, 2, 'neigh_op_tnr_4')
// (7, 2, 'sp4_r_v_b_37')
// (7, 3, 'neigh_op_rgt_4')
// (7, 3, 'sp4_r_v_b_24')
// (7, 4, 'neigh_op_bnr_4')
// (7, 4, 'sp4_r_v_b_13')
// (7, 5, 'sp4_r_v_b_0')
// (8, 1, 'sp4_v_t_37')
// (8, 2, 'neigh_op_top_4')
// (8, 2, 'sp4_v_b_37')
// (8, 3, 'lutff_4/out')
// (8, 3, 'sp4_v_b_24')
// (8, 4, 'local_g0_4')
// (8, 4, 'lutff_0/in_2')
// (8, 4, 'neigh_op_bot_4')
// (8, 4, 'sp4_v_b_13')
// (8, 5, 'local_g1_0')
// (8, 5, 'lutff_2/in_1')
// (8, 5, 'sp4_v_b_0')
// (9, 2, 'neigh_op_tnl_4')
// (9, 3, 'neigh_op_lft_4')
// (9, 4, 'neigh_op_bnl_4')

wire n415;
// (7, 2, 'neigh_op_tnr_6')
// (7, 3, 'neigh_op_rgt_6')
// (7, 4, 'neigh_op_bnr_6')
// (8, 2, 'neigh_op_top_6')
// (8, 3, 'local_g3_6')
// (8, 3, 'lutff_4/in_3')
// (8, 3, 'lutff_6/out')
// (8, 4, 'neigh_op_bot_6')
// (9, 2, 'neigh_op_tnl_6')
// (9, 3, 'neigh_op_lft_6')
// (9, 4, 'neigh_op_bnl_6')

wire n416;
// (7, 2, 'sp4_r_v_b_44')
// (7, 3, 'sp4_r_v_b_33')
// (7, 4, 'sp4_r_v_b_20')
// (7, 5, 'sp4_r_v_b_9')
// (8, 1, 'sp4_v_t_44')
// (8, 2, 'sp4_v_b_44')
// (8, 3, 'local_g3_1')
// (8, 3, 'lutff_5/in_3')
// (8, 3, 'lutff_7/in_3')
// (8, 3, 'sp4_v_b_33')
// (8, 4, 'neigh_op_tnr_2')
// (8, 4, 'sp4_v_b_20')
// (8, 5, 'neigh_op_rgt_2')
// (8, 5, 'sp4_h_r_9')
// (8, 5, 'sp4_v_b_9')
// (8, 6, 'neigh_op_bnr_2')
// (9, 4, 'neigh_op_top_2')
// (9, 5, 'lutff_2/out')
// (9, 5, 'sp4_h_r_20')
// (9, 6, 'neigh_op_bot_2')
// (10, 4, 'neigh_op_tnl_2')
// (10, 5, 'neigh_op_lft_2')
// (10, 5, 'sp4_h_r_33')
// (10, 6, 'neigh_op_bnl_2')
// (11, 5, 'sp4_h_r_44')
// (12, 5, 'sp4_h_l_44')

wire n417;
// (7, 3, 'neigh_op_tnr_0')
// (7, 4, 'neigh_op_rgt_0')
// (7, 5, 'neigh_op_bnr_0')
// (8, 3, 'neigh_op_top_0')
// (8, 4, 'local_g0_0')
// (8, 4, 'lutff_0/out')
// (8, 4, 'lutff_7/in_1')
// (8, 5, 'neigh_op_bot_0')
// (9, 3, 'neigh_op_tnl_0')
// (9, 4, 'neigh_op_lft_0')
// (9, 5, 'neigh_op_bnl_0')

wire n418;
// (7, 3, 'neigh_op_tnr_2')
// (7, 4, 'neigh_op_rgt_2')
// (7, 5, 'neigh_op_bnr_2')
// (8, 3, 'local_g0_2')
// (8, 3, 'local_g1_2')
// (8, 3, 'lutff_3/in_2')
// (8, 3, 'lutff_7/in_1')
// (8, 3, 'neigh_op_top_2')
// (8, 4, 'local_g1_2')
// (8, 4, 'lutff_2/out')
// (8, 4, 'lutff_3/in_2')
// (8, 5, 'neigh_op_bot_2')
// (9, 3, 'local_g2_2')
// (9, 3, 'lutff_7/in_1')
// (9, 3, 'neigh_op_tnl_2')
// (9, 4, 'neigh_op_lft_2')
// (9, 5, 'neigh_op_bnl_2')

wire n419;
// (7, 3, 'neigh_op_tnr_4')
// (7, 4, 'local_g2_4')
// (7, 4, 'local_g3_4')
// (7, 4, 'lutff_0/in_3')
// (7, 4, 'lutff_5/in_1')
// (7, 4, 'neigh_op_rgt_4')
// (7, 5, 'neigh_op_bnr_4')
// (8, 3, 'local_g0_4')
// (8, 3, 'local_g1_4')
// (8, 3, 'lutff_1/in_1')
// (8, 3, 'lutff_2/in_3')
// (8, 3, 'neigh_op_top_4')
// (8, 4, 'lutff_4/out')
// (8, 5, 'neigh_op_bot_4')
// (9, 3, 'neigh_op_tnl_4')
// (9, 4, 'neigh_op_lft_4')
// (9, 5, 'neigh_op_bnl_4')

wire n420;
// (7, 3, 'neigh_op_tnr_6')
// (7, 4, 'neigh_op_rgt_6')
// (7, 5, 'neigh_op_bnr_6')
// (8, 3, 'neigh_op_top_6')
// (8, 4, 'local_g0_6')
// (8, 4, 'local_g1_6')
// (8, 4, 'lutff_1/in_1')
// (8, 4, 'lutff_4/in_1')
// (8, 4, 'lutff_6/out')
// (8, 5, 'neigh_op_bot_6')
// (9, 3, 'neigh_op_tnl_6')
// (9, 4, 'local_g0_6')
// (9, 4, 'lutff_6/in_0')
// (9, 4, 'neigh_op_lft_6')
// (9, 5, 'neigh_op_bnl_6')

wire n421;
// (7, 4, 'neigh_op_tnr_0')
// (7, 5, 'neigh_op_rgt_0')
// (7, 6, 'neigh_op_bnr_0')
// (8, 2, 'sp4_r_v_b_36')
// (8, 3, 'sp4_r_v_b_25')
// (8, 4, 'neigh_op_top_0')
// (8, 4, 'sp4_r_v_b_12')
// (8, 5, 'lutff_0/out')
// (8, 5, 'sp4_h_r_0')
// (8, 5, 'sp4_r_v_b_1')
// (8, 6, 'neigh_op_bot_0')
// (8, 6, 'sp4_r_v_b_36')
// (8, 7, 'sp4_r_v_b_25')
// (8, 8, 'sp4_r_v_b_12')
// (8, 9, 'sp4_r_v_b_1')
// (8, 10, 'sp4_r_v_b_36')
// (8, 11, 'sp4_r_v_b_25')
// (8, 12, 'sp4_r_v_b_12')
// (8, 13, 'sp4_r_v_b_1')
// (9, 1, 'sp4_v_t_36')
// (9, 2, 'sp4_v_b_36')
// (9, 3, 'sp4_v_b_25')
// (9, 4, 'neigh_op_tnl_0')
// (9, 4, 'sp4_v_b_12')
// (9, 5, 'neigh_op_lft_0')
// (9, 5, 'sp4_h_r_13')
// (9, 5, 'sp4_v_b_1')
// (9, 5, 'sp4_v_t_36')
// (9, 6, 'neigh_op_bnl_0')
// (9, 6, 'sp4_v_b_36')
// (9, 7, 'sp4_v_b_25')
// (9, 8, 'sp4_v_b_12')
// (9, 9, 'local_g0_1')
// (9, 9, 'lutff_5/in_2')
// (9, 9, 'sp4_v_b_1')
// (9, 9, 'sp4_v_t_36')
// (9, 10, 'sp4_v_b_36')
// (9, 11, 'sp4_v_b_25')
// (9, 12, 'sp4_v_b_12')
// (9, 13, 'local_g0_1')
// (9, 13, 'lutff_5/in_0')
// (9, 13, 'sp4_v_b_1')
// (10, 5, 'sp4_h_r_24')
// (11, 5, 'sp4_h_r_37')
// (11, 6, 'sp4_r_v_b_40')
// (11, 7, 'sp4_r_v_b_29')
// (11, 8, 'sp4_r_v_b_16')
// (11, 9, 'sp4_r_v_b_5')
// (11, 10, 'sp4_r_v_b_36')
// (11, 11, 'local_g0_1')
// (11, 11, 'lutff_3/in_2')
// (11, 11, 'lutff_7/in_2')
// (11, 11, 'sp4_r_v_b_25')
// (11, 12, 'sp4_r_v_b_12')
// (11, 13, 'sp4_r_v_b_1')
// (12, 5, 'sp4_h_l_37')
// (12, 5, 'sp4_v_t_40')
// (12, 6, 'sp4_v_b_40')
// (12, 7, 'sp4_v_b_29')
// (12, 8, 'sp4_v_b_16')
// (12, 9, 'sp4_v_b_5')
// (12, 9, 'sp4_v_t_36')
// (12, 10, 'sp4_v_b_36')
// (12, 11, 'sp4_v_b_25')
// (12, 12, 'sp4_v_b_12')
// (12, 13, 'sp4_v_b_1')

wire n422;
// (7, 4, 'neigh_op_tnr_1')
// (7, 5, 'neigh_op_rgt_1')
// (7, 6, 'neigh_op_bnr_1')
// (8, 4, 'neigh_op_top_1')
// (8, 5, 'local_g1_1')
// (8, 5, 'lutff_1/out')
// (8, 5, 'lutff_3/in_1')
// (8, 6, 'neigh_op_bot_1')
// (9, 4, 'neigh_op_tnl_1')
// (9, 5, 'neigh_op_lft_1')
// (9, 6, 'neigh_op_bnl_1')

wire n423;
// (7, 4, 'neigh_op_tnr_2')
// (7, 5, 'neigh_op_rgt_2')
// (7, 5, 'sp4_r_v_b_36')
// (7, 6, 'neigh_op_bnr_2')
// (7, 6, 'sp4_r_v_b_25')
// (7, 7, 'sp4_r_v_b_12')
// (7, 8, 'sp4_r_v_b_1')
// (8, 4, 'neigh_op_top_2')
// (8, 4, 'sp4_v_t_36')
// (8, 5, 'lutff_2/out')
// (8, 5, 'sp4_r_v_b_37')
// (8, 5, 'sp4_v_b_36')
// (8, 6, 'neigh_op_bot_2')
// (8, 6, 'sp4_r_v_b_24')
// (8, 6, 'sp4_v_b_25')
// (8, 7, 'local_g0_4')
// (8, 7, 'lutff_0/in_2')
// (8, 7, 'sp4_r_v_b_13')
// (8, 7, 'sp4_v_b_12')
// (8, 8, 'sp4_h_r_1')
// (8, 8, 'sp4_r_v_b_0')
// (8, 8, 'sp4_v_b_1')
// (9, 4, 'neigh_op_tnl_2')
// (9, 4, 'sp4_v_t_37')
// (9, 5, 'neigh_op_lft_2')
// (9, 5, 'sp4_v_b_37')
// (9, 6, 'neigh_op_bnl_2')
// (9, 6, 'sp4_v_b_24')
// (9, 7, 'sp4_v_b_13')
// (9, 8, 'local_g1_0')
// (9, 8, 'lutff_3/in_0')
// (9, 8, 'sp4_h_r_12')
// (9, 8, 'sp4_v_b_0')
// (10, 8, 'sp4_h_r_25')
// (11, 8, 'sp4_h_r_36')
// (11, 9, 'sp4_r_v_b_36')
// (11, 10, 'local_g0_1')
// (11, 10, 'local_g1_1')
// (11, 10, 'lutff_1/in_2')
// (11, 10, 'lutff_2/in_2')
// (11, 10, 'sp4_r_v_b_25')
// (11, 11, 'sp4_r_v_b_12')
// (11, 12, 'sp4_r_v_b_1')
// (12, 8, 'sp4_h_l_36')
// (12, 8, 'sp4_v_t_36')
// (12, 9, 'sp4_v_b_36')
// (12, 10, 'sp4_v_b_25')
// (12, 11, 'sp4_v_b_12')
// (12, 12, 'sp4_v_b_1')

wire n424;
// (7, 4, 'neigh_op_tnr_3')
// (7, 5, 'neigh_op_rgt_3')
// (7, 6, 'neigh_op_bnr_3')
// (8, 0, 'span12_vert_14')
// (8, 1, 'sp12_v_b_14')
// (8, 2, 'sp12_v_b_13')
// (8, 3, 'local_g2_2')
// (8, 3, 'local_g3_2')
// (8, 3, 'lutff_3/in_3')
// (8, 3, 'lutff_5/in_2')
// (8, 3, 'sp12_v_b_10')
// (8, 4, 'neigh_op_top_3')
// (8, 4, 'sp12_v_b_9')
// (8, 5, 'lutff_3/out')
// (8, 5, 'sp12_v_b_6')
// (8, 6, 'neigh_op_bot_3')
// (8, 6, 'sp12_v_b_5')
// (8, 7, 'sp12_v_b_2')
// (8, 8, 'sp12_v_b_1')
// (9, 4, 'local_g3_3')
// (9, 4, 'lutff_6/in_2')
// (9, 4, 'neigh_op_tnl_3')
// (9, 5, 'neigh_op_lft_3')
// (9, 6, 'neigh_op_bnl_3')

wire n425;
// (7, 4, 'neigh_op_tnr_4')
// (7, 5, 'neigh_op_rgt_4')
// (7, 6, 'neigh_op_bnr_4')
// (8, 4, 'neigh_op_top_4')
// (8, 5, 'local_g1_4')
// (8, 5, 'lutff_3/in_0')
// (8, 5, 'lutff_4/out')
// (8, 5, 'lutff_5/in_2')
// (8, 6, 'neigh_op_bot_4')
// (9, 4, 'neigh_op_tnl_4')
// (9, 5, 'neigh_op_lft_4')
// (9, 6, 'neigh_op_bnl_4')

wire n426;
// (7, 4, 'neigh_op_tnr_6')
// (7, 5, 'neigh_op_rgt_6')
// (7, 6, 'neigh_op_bnr_6')
// (8, 4, 'neigh_op_top_6')
// (8, 5, 'lutff_6/out')
// (8, 6, 'neigh_op_bot_6')
// (9, 4, 'neigh_op_tnl_6')
// (9, 5, 'local_g0_6')
// (9, 5, 'local_g1_6')
// (9, 5, 'lutff_3/in_3')
// (9, 5, 'lutff_6/in_3')
// (9, 5, 'neigh_op_lft_6')
// (9, 6, 'neigh_op_bnl_6')

reg n427 = 0;
// (7, 4, 'neigh_op_tnr_7')
// (7, 5, 'neigh_op_rgt_7')
// (7, 6, 'neigh_op_bnr_7')
// (8, 4, 'neigh_op_top_7')
// (8, 5, 'lutff_7/out')
// (8, 6, 'local_g1_7')
// (8, 6, 'lutff_6/in_0')
// (8, 6, 'neigh_op_bot_7')
// (9, 4, 'neigh_op_tnl_7')
// (9, 5, 'neigh_op_lft_7')
// (9, 6, 'neigh_op_bnl_7')

reg n428 = 0;
// (7, 4, 'sp4_r_v_b_40')
// (7, 5, 'neigh_op_tnr_0')
// (7, 5, 'sp4_r_v_b_29')
// (7, 6, 'local_g2_0')
// (7, 6, 'lutff_6/in_0')
// (7, 6, 'neigh_op_rgt_0')
// (7, 6, 'sp4_r_v_b_16')
// (7, 7, 'neigh_op_bnr_0')
// (7, 7, 'sp4_r_v_b_5')
// (7, 8, 'sp4_r_v_b_36')
// (7, 9, 'local_g0_1')
// (7, 9, 'lutff_1/in_2')
// (7, 9, 'lutff_7/in_2')
// (7, 9, 'sp4_r_v_b_25')
// (7, 10, 'sp4_r_v_b_12')
// (7, 11, 'sp4_r_v_b_1')
// (8, 2, 'sp12_v_t_23')
// (8, 3, 'sp12_v_b_23')
// (8, 3, 'sp4_v_t_40')
// (8, 4, 'sp12_v_b_20')
// (8, 4, 'sp4_v_b_40')
// (8, 5, 'neigh_op_top_0')
// (8, 5, 'sp12_v_b_19')
// (8, 5, 'sp4_v_b_29')
// (8, 6, 'lutff_0/out')
// (8, 6, 'sp12_v_b_16')
// (8, 6, 'sp4_v_b_16')
// (8, 7, 'neigh_op_bot_0')
// (8, 7, 'sp12_v_b_15')
// (8, 7, 'sp4_v_b_5')
// (8, 7, 'sp4_v_t_36')
// (8, 8, 'sp12_v_b_12')
// (8, 8, 'sp4_v_b_36')
// (8, 9, 'local_g3_3')
// (8, 9, 'lutff_4/in_0')
// (8, 9, 'sp12_v_b_11')
// (8, 9, 'sp4_v_b_25')
// (8, 10, 'sp12_v_b_8')
// (8, 10, 'sp4_v_b_12')
// (8, 11, 'sp12_v_b_7')
// (8, 11, 'sp4_v_b_1')
// (8, 12, 'sp12_v_b_4')
// (8, 13, 'sp12_v_b_3')
// (8, 14, 'sp12_v_b_0')
// (9, 5, 'neigh_op_tnl_0')
// (9, 6, 'neigh_op_lft_0')
// (9, 7, 'neigh_op_bnl_0')

reg n429 = 0;
// (7, 4, 'sp4_r_v_b_41')
// (7, 5, 'sp4_r_v_b_28')
// (7, 6, 'neigh_op_tnr_2')
// (7, 6, 'sp4_r_v_b_17')
// (7, 7, 'neigh_op_rgt_2')
// (7, 7, 'sp4_r_v_b_4')
// (7, 8, 'neigh_op_bnr_2')
// (8, 3, 'sp4_v_t_41')
// (8, 4, 'sp4_v_b_41')
// (8, 5, 'local_g3_4')
// (8, 5, 'lutff_0/in_3')
// (8, 5, 'sp4_v_b_28')
// (8, 6, 'neigh_op_top_2')
// (8, 6, 'sp4_v_b_17')
// (8, 7, 'lutff_2/out')
// (8, 7, 'sp4_v_b_4')
// (8, 8, 'neigh_op_bot_2')
// (9, 6, 'neigh_op_tnl_2')
// (9, 7, 'neigh_op_lft_2')
// (9, 8, 'neigh_op_bnl_2')

reg n430 = 0;
// (7, 4, 'sp4_r_v_b_45')
// (7, 5, 'sp4_r_v_b_32')
// (7, 6, 'neigh_op_tnr_4')
// (7, 6, 'sp4_r_v_b_21')
// (7, 7, 'neigh_op_rgt_4')
// (7, 7, 'sp4_r_v_b_8')
// (7, 8, 'neigh_op_bnr_4')
// (8, 3, 'sp4_v_t_45')
// (8, 4, 'sp4_v_b_45')
// (8, 5, 'local_g3_0')
// (8, 5, 'lutff_2/in_3')
// (8, 5, 'sp4_v_b_32')
// (8, 6, 'neigh_op_top_4')
// (8, 6, 'sp4_v_b_21')
// (8, 7, 'lutff_4/out')
// (8, 7, 'sp4_v_b_8')
// (8, 8, 'neigh_op_bot_4')
// (9, 6, 'neigh_op_tnl_4')
// (9, 7, 'neigh_op_lft_4')
// (9, 8, 'neigh_op_bnl_4')

reg n431 = 0;
// (7, 5, 'local_g3_7')
// (7, 5, 'lutff_5/in_3')
// (7, 5, 'neigh_op_tnr_7')
// (7, 6, 'neigh_op_rgt_7')
// (7, 7, 'neigh_op_bnr_7')
// (8, 5, 'neigh_op_top_7')
// (8, 6, 'lutff_7/out')
// (8, 7, 'neigh_op_bot_7')
// (9, 5, 'neigh_op_tnl_7')
// (9, 6, 'neigh_op_lft_7')
// (9, 7, 'neigh_op_bnl_7')

reg n432 = 0;
// (7, 5, 'neigh_op_tnr_1')
// (7, 6, 'neigh_op_rgt_1')
// (7, 7, 'neigh_op_bnr_1')
// (8, 5, 'neigh_op_top_1')
// (8, 6, 'local_g0_1')
// (8, 6, 'lutff_1/out')
// (8, 6, 'lutff_7/in_0')
// (8, 7, 'neigh_op_bot_1')
// (9, 5, 'neigh_op_tnl_1')
// (9, 6, 'neigh_op_lft_1')
// (9, 7, 'neigh_op_bnl_1')

reg n433 = 0;
// (7, 5, 'neigh_op_tnr_3')
// (7, 6, 'neigh_op_rgt_3')
// (7, 7, 'neigh_op_bnr_3')
// (8, 5, 'neigh_op_top_3')
// (8, 6, 'local_g0_3')
// (8, 6, 'lutff_3/out')
// (8, 6, 'lutff_5/in_0')
// (8, 7, 'neigh_op_bot_3')
// (9, 5, 'neigh_op_tnl_3')
// (9, 6, 'neigh_op_lft_3')
// (9, 7, 'neigh_op_bnl_3')

reg n434 = 0;
// (7, 5, 'neigh_op_tnr_4')
// (7, 6, 'neigh_op_rgt_4')
// (7, 7, 'neigh_op_bnr_4')
// (8, 0, 'span12_vert_19')
// (8, 1, 'sp12_v_b_19')
// (8, 2, 'sp12_v_b_16')
// (8, 3, 'sp12_v_b_15')
// (8, 4, 'sp12_v_b_12')
// (8, 5, 'local_g2_3')
// (8, 5, 'lutff_4/in_3')
// (8, 5, 'neigh_op_top_4')
// (8, 5, 'sp12_v_b_11')
// (8, 6, 'local_g0_4')
// (8, 6, 'lutff_2/in_0')
// (8, 6, 'lutff_4/out')
// (8, 6, 'sp12_v_b_8')
// (8, 7, 'neigh_op_bot_4')
// (8, 7, 'sp12_v_b_7')
// (8, 8, 'sp12_v_b_4')
// (8, 9, 'sp12_v_b_3')
// (8, 10, 'sp12_v_b_0')
// (9, 5, 'neigh_op_tnl_4')
// (9, 6, 'neigh_op_lft_4')
// (9, 7, 'neigh_op_bnl_4')

reg n435 = 0;
// (7, 5, 'neigh_op_tnr_5')
// (7, 6, 'neigh_op_rgt_5')
// (7, 7, 'neigh_op_bnr_5')
// (8, 5, 'neigh_op_top_5')
// (8, 6, 'local_g0_5')
// (8, 6, 'lutff_1/in_0')
// (8, 6, 'lutff_5/out')
// (8, 7, 'neigh_op_bot_5')
// (9, 5, 'neigh_op_tnl_5')
// (9, 6, 'neigh_op_lft_5')
// (9, 7, 'neigh_op_bnl_5')

reg n436 = 0;
// (7, 5, 'neigh_op_tnr_6')
// (7, 6, 'neigh_op_rgt_6')
// (7, 7, 'neigh_op_bnr_6')
// (8, 5, 'neigh_op_top_6')
// (8, 6, 'local_g2_6')
// (8, 6, 'lutff_4/in_0')
// (8, 6, 'lutff_6/out')
// (8, 7, 'neigh_op_bot_6')
// (9, 5, 'neigh_op_tnl_6')
// (9, 6, 'neigh_op_lft_6')
// (9, 7, 'neigh_op_bnl_6')

wire n437;
// (7, 5, 'sp4_h_r_7')
// (8, 5, 'local_g0_2')
// (8, 5, 'lutff_3/in_3')
// (8, 5, 'lutff_5/in_3')
// (8, 5, 'sp4_h_r_18')
// (9, 5, 'sp4_h_r_31')
// (10, 2, 'sp4_r_v_b_39')
// (10, 3, 'sp4_r_v_b_26')
// (10, 4, 'neigh_op_tnr_1')
// (10, 4, 'sp4_r_v_b_15')
// (10, 5, 'neigh_op_rgt_1')
// (10, 5, 'sp4_h_r_42')
// (10, 5, 'sp4_r_v_b_2')
// (10, 6, 'neigh_op_bnr_1')
// (11, 1, 'sp4_v_t_39')
// (11, 2, 'sp4_v_b_39')
// (11, 3, 'sp4_v_b_26')
// (11, 4, 'neigh_op_top_1')
// (11, 4, 'sp4_v_b_15')
// (11, 5, 'lutff_1/out')
// (11, 5, 'sp4_h_l_42')
// (11, 5, 'sp4_v_b_2')
// (11, 6, 'neigh_op_bot_1')
// (12, 4, 'neigh_op_tnl_1')
// (12, 5, 'neigh_op_lft_1')
// (12, 6, 'neigh_op_bnl_1')

reg n438 = 0;
// (7, 6, 'neigh_op_tnr_0')
// (7, 7, 'neigh_op_rgt_0')
// (7, 8, 'neigh_op_bnr_0')
// (8, 6, 'neigh_op_top_0')
// (8, 7, 'local_g0_0')
// (8, 7, 'lutff_0/out')
// (8, 7, 'lutff_6/in_0')
// (8, 8, 'neigh_op_bot_0')
// (9, 6, 'neigh_op_tnl_0')
// (9, 7, 'neigh_op_lft_0')
// (9, 8, 'neigh_op_bnl_0')

reg n439 = 0;
// (7, 6, 'neigh_op_tnr_1')
// (7, 7, 'neigh_op_rgt_1')
// (7, 8, 'neigh_op_bnr_1')
// (8, 6, 'neigh_op_top_1')
// (8, 7, 'local_g1_1')
// (8, 7, 'lutff_1/out')
// (8, 7, 'lutff_4/in_0')
// (8, 8, 'neigh_op_bot_1')
// (9, 6, 'neigh_op_tnl_1')
// (9, 7, 'neigh_op_lft_1')
// (9, 8, 'neigh_op_bnl_1')

reg n440 = 0;
// (7, 6, 'neigh_op_tnr_3')
// (7, 7, 'local_g2_3')
// (7, 7, 'lutff_0/in_3')
// (7, 7, 'neigh_op_rgt_3')
// (7, 8, 'neigh_op_bnr_3')
// (8, 6, 'neigh_op_top_3')
// (8, 7, 'lutff_3/out')
// (8, 8, 'neigh_op_bot_3')
// (9, 6, 'neigh_op_tnl_3')
// (9, 7, 'neigh_op_lft_3')
// (9, 8, 'neigh_op_bnl_3')

reg n441 = 0;
// (7, 6, 'neigh_op_tnr_5')
// (7, 7, 'neigh_op_rgt_5')
// (7, 8, 'neigh_op_bnr_5')
// (8, 6, 'neigh_op_top_5')
// (8, 7, 'local_g1_5')
// (8, 7, 'lutff_2/in_0')
// (8, 7, 'lutff_5/out')
// (8, 8, 'neigh_op_bot_5')
// (9, 6, 'neigh_op_tnl_5')
// (9, 7, 'neigh_op_lft_5')
// (9, 8, 'neigh_op_bnl_5')

reg n442 = 0;
// (7, 6, 'neigh_op_tnr_6')
// (7, 7, 'neigh_op_rgt_6')
// (7, 8, 'neigh_op_bnr_6')
// (8, 6, 'neigh_op_top_6')
// (8, 7, 'local_g1_6')
// (8, 7, 'lutff_1/in_0')
// (8, 7, 'lutff_6/out')
// (8, 8, 'neigh_op_bot_6')
// (9, 6, 'neigh_op_tnl_6')
// (9, 7, 'neigh_op_lft_6')
// (9, 8, 'neigh_op_bnl_6')

reg n443 = 0;
// (7, 6, 'neigh_op_tnr_7')
// (7, 7, 'neigh_op_rgt_7')
// (7, 8, 'neigh_op_bnr_7')
// (8, 6, 'neigh_op_top_7')
// (8, 7, 'local_g0_7')
// (8, 7, 'lutff_3/in_0')
// (8, 7, 'lutff_7/out')
// (8, 8, 'neigh_op_bot_7')
// (9, 6, 'neigh_op_tnl_7')
// (9, 7, 'neigh_op_lft_7')
// (9, 8, 'neigh_op_bnl_7')

reg n444 = 0;
// (7, 6, 'sp4_h_r_10')
// (8, 5, 'neigh_op_tnr_1')
// (8, 6, 'neigh_op_rgt_1')
// (8, 6, 'sp4_h_r_23')
// (8, 7, 'neigh_op_bnr_1')
// (9, 5, 'neigh_op_top_1')
// (9, 6, 'lutff_1/out')
// (9, 6, 'sp4_h_r_34')
// (9, 7, 'neigh_op_bot_1')
// (10, 3, 'sp4_r_v_b_41')
// (10, 4, 'sp4_r_v_b_28')
// (10, 5, 'neigh_op_tnl_1')
// (10, 5, 'sp4_r_v_b_17')
// (10, 6, 'neigh_op_lft_1')
// (10, 6, 'sp4_h_r_47')
// (10, 6, 'sp4_r_v_b_4')
// (10, 7, 'neigh_op_bnl_1')
// (11, 2, 'sp4_v_t_41')
// (11, 3, 'sp4_v_b_41')
// (11, 4, 'sp4_v_b_28')
// (11, 5, 'local_g0_1')
// (11, 5, 'lutff_5/in_0')
// (11, 5, 'sp4_v_b_17')
// (11, 6, 'sp4_h_l_47')
// (11, 6, 'sp4_v_b_4')

reg n445 = 0;
// (7, 6, 'sp4_h_r_4')
// (8, 6, 'local_g1_1')
// (8, 6, 'lutff_3/in_3')
// (8, 6, 'sp4_h_r_17')
// (9, 6, 'sp4_h_r_28')
// (10, 6, 'sp4_h_r_41')
// (11, 5, 'neigh_op_tnr_6')
// (11, 6, 'neigh_op_rgt_6')
// (11, 6, 'sp4_h_l_41')
// (11, 6, 'sp4_h_r_1')
// (11, 7, 'neigh_op_bnr_6')
// (12, 5, 'neigh_op_top_6')
// (12, 6, 'lutff_6/out')
// (12, 6, 'sp4_h_r_12')
// (12, 7, 'neigh_op_bot_6')
// (13, 5, 'logic_op_tnl_6')
// (13, 6, 'logic_op_lft_6')
// (13, 6, 'span4_horz_12')
// (13, 7, 'logic_op_bnl_6')

wire n446;
// (7, 7, 'neigh_op_tnr_0')
// (7, 8, 'neigh_op_rgt_0')
// (7, 9, 'neigh_op_bnr_0')
// (8, 5, 'sp4_r_v_b_36')
// (8, 6, 'sp4_r_v_b_25')
// (8, 7, 'neigh_op_top_0')
// (8, 7, 'sp4_r_v_b_12')
// (8, 8, 'local_g1_0')
// (8, 8, 'lutff_0/out')
// (8, 8, 'lutff_5/in_2')
// (8, 8, 'lutff_7/in_2')
// (8, 8, 'sp4_r_v_b_1')
// (8, 9, 'neigh_op_bot_0')
// (9, 4, 'sp4_v_t_36')
// (9, 5, 'sp4_v_b_36')
// (9, 6, 'sp4_v_b_25')
// (9, 7, 'neigh_op_tnl_0')
// (9, 7, 'sp4_v_b_12')
// (9, 8, 'local_g0_0')
// (9, 8, 'local_g0_1')
// (9, 8, 'lutff_1/in_2')
// (9, 8, 'lutff_6/in_0')
// (9, 8, 'neigh_op_lft_0')
// (9, 8, 'sp4_v_b_1')
// (9, 9, 'neigh_op_bnl_0')

reg n447 = 0;
// (7, 7, 'neigh_op_tnr_1')
// (7, 8, 'neigh_op_rgt_1')
// (7, 9, 'neigh_op_bnr_1')
// (8, 5, 'sp4_r_v_b_38')
// (8, 6, 'sp4_r_v_b_27')
// (8, 7, 'neigh_op_top_1')
// (8, 7, 'sp4_r_v_b_14')
// (8, 8, 'local_g1_3')
// (8, 8, 'lutff_1/out')
// (8, 8, 'lutff_2/in_0')
// (8, 8, 'sp4_r_v_b_3')
// (8, 9, 'neigh_op_bot_1')
// (9, 4, 'sp4_v_t_38')
// (9, 5, 'sp4_v_b_38')
// (9, 6, 'sp4_v_b_27')
// (9, 7, 'neigh_op_tnl_1')
// (9, 7, 'sp4_v_b_14')
// (9, 8, 'neigh_op_lft_1')
// (9, 8, 'sp4_v_b_3')
// (9, 9, 'neigh_op_bnl_1')

reg n448 = 0;
// (7, 7, 'neigh_op_tnr_2')
// (7, 8, 'neigh_op_rgt_2')
// (7, 9, 'neigh_op_bnr_2')
// (8, 7, 'neigh_op_top_2')
// (8, 8, 'local_g0_2')
// (8, 8, 'lutff_2/out')
// (8, 8, 'lutff_6/in_0')
// (8, 9, 'neigh_op_bot_2')
// (9, 7, 'neigh_op_tnl_2')
// (9, 8, 'neigh_op_lft_2')
// (9, 9, 'neigh_op_bnl_2')

reg n449 = 0;
// (7, 7, 'neigh_op_tnr_5')
// (7, 8, 'neigh_op_rgt_5')
// (7, 9, 'neigh_op_bnr_5')
// (8, 7, 'neigh_op_top_5')
// (8, 8, 'local_g0_5')
// (8, 8, 'lutff_1/in_0')
// (8, 8, 'lutff_5/out')
// (8, 9, 'neigh_op_bot_5')
// (9, 7, 'neigh_op_tnl_5')
// (9, 8, 'neigh_op_lft_5')
// (9, 9, 'neigh_op_bnl_5')

reg n450 = 0;
// (7, 7, 'neigh_op_tnr_6')
// (7, 8, 'neigh_op_rgt_6')
// (7, 9, 'neigh_op_bnr_6')
// (8, 7, 'neigh_op_top_6')
// (8, 8, 'local_g1_6')
// (8, 8, 'lutff_0/in_3')
// (8, 8, 'lutff_6/out')
// (8, 9, 'neigh_op_bot_6')
// (9, 7, 'neigh_op_tnl_6')
// (9, 8, 'neigh_op_lft_6')
// (9, 9, 'neigh_op_bnl_6')

reg n451 = 0;
// (7, 7, 'neigh_op_tnr_7')
// (7, 8, 'neigh_op_rgt_7')
// (7, 9, 'neigh_op_bnr_7')
// (8, 7, 'neigh_op_top_7')
// (8, 8, 'lutff_7/out')
// (8, 9, 'neigh_op_bot_7')
// (9, 7, 'neigh_op_tnl_7')
// (9, 8, 'local_g1_7')
// (9, 8, 'lutff_1/in_1')
// (9, 8, 'neigh_op_lft_7')
// (9, 9, 'neigh_op_bnl_7')

wire n452;
// (7, 8, 'neigh_op_tnr_0')
// (7, 9, 'local_g2_0')
// (7, 9, 'lutff_1/in_3')
// (7, 9, 'neigh_op_rgt_0')
// (7, 10, 'neigh_op_bnr_0')
// (8, 8, 'neigh_op_top_0')
// (8, 9, 'lutff_0/out')
// (8, 10, 'neigh_op_bot_0')
// (9, 8, 'neigh_op_tnl_0')
// (9, 9, 'neigh_op_lft_0')
// (9, 10, 'neigh_op_bnl_0')

wire n453;
// (7, 8, 'neigh_op_tnr_1')
// (7, 9, 'neigh_op_rgt_1')
// (7, 10, 'neigh_op_bnr_1')
// (8, 8, 'neigh_op_top_1')
// (8, 9, 'local_g2_1')
// (8, 9, 'lutff_0/in_3')
// (8, 9, 'lutff_1/out')
// (8, 10, 'neigh_op_bot_1')
// (9, 8, 'neigh_op_tnl_1')
// (9, 9, 'neigh_op_lft_1')
// (9, 10, 'neigh_op_bnl_1')

reg n454 = 0;
// (7, 8, 'neigh_op_tnr_2')
// (7, 9, 'neigh_op_rgt_2')
// (7, 9, 'sp4_h_r_9')
// (7, 10, 'neigh_op_bnr_2')
// (8, 8, 'neigh_op_top_2')
// (8, 9, 'lutff_2/out')
// (8, 9, 'sp4_h_r_20')
// (8, 10, 'neigh_op_bot_2')
// (9, 8, 'neigh_op_tnl_2')
// (9, 9, 'neigh_op_lft_2')
// (9, 9, 'sp4_h_r_33')
// (9, 10, 'neigh_op_bnl_2')
// (10, 6, 'sp4_r_v_b_44')
// (10, 7, 'sp4_r_v_b_33')
// (10, 8, 'sp4_r_v_b_20')
// (10, 9, 'sp4_h_r_44')
// (10, 9, 'sp4_r_v_b_9')
// (11, 5, 'sp4_v_t_44')
// (11, 6, 'sp4_v_b_44')
// (11, 7, 'sp4_v_b_33')
// (11, 8, 'local_g1_4')
// (11, 8, 'lutff_3/in_0')
// (11, 8, 'sp4_v_b_20')
// (11, 9, 'sp4_h_l_44')
// (11, 9, 'sp4_v_b_9')

reg n455 = 0;
// (7, 8, 'neigh_op_tnr_3')
// (7, 9, 'neigh_op_rgt_3')
// (7, 10, 'neigh_op_bnr_3')
// (8, 8, 'neigh_op_top_3')
// (8, 9, 'lutff_3/out')
// (8, 10, 'neigh_op_bot_3')
// (9, 8, 'neigh_op_tnl_3')
// (9, 9, 'local_g1_3')
// (9, 9, 'lutff_4/in_0')
// (9, 9, 'neigh_op_lft_3')
// (9, 10, 'neigh_op_bnl_3')

reg n456 = 0;
// (7, 8, 'neigh_op_tnr_4')
// (7, 9, 'neigh_op_rgt_4')
// (7, 10, 'neigh_op_bnr_4')
// (8, 8, 'neigh_op_top_4')
// (8, 9, 'lutff_4/out')
// (8, 9, 'sp4_h_r_8')
// (8, 10, 'neigh_op_bot_4')
// (9, 8, 'neigh_op_tnl_4')
// (9, 9, 'neigh_op_lft_4')
// (9, 9, 'sp4_h_r_21')
// (9, 10, 'neigh_op_bnl_4')
// (10, 9, 'sp4_h_r_32')
// (11, 9, 'local_g2_5')
// (11, 9, 'lutff_3/in_0')
// (11, 9, 'sp4_h_r_45')
// (12, 9, 'sp4_h_l_45')

reg n457 = 0;
// (7, 8, 'neigh_op_tnr_6')
// (7, 9, 'neigh_op_rgt_6')
// (7, 10, 'neigh_op_bnr_6')
// (8, 8, 'neigh_op_top_6')
// (8, 9, 'local_g2_6')
// (8, 9, 'lutff_2/in_0')
// (8, 9, 'lutff_6/out')
// (8, 10, 'neigh_op_bot_6')
// (9, 8, 'neigh_op_tnl_6')
// (9, 9, 'neigh_op_lft_6')
// (9, 10, 'neigh_op_bnl_6')

reg n458 = 0;
// (7, 8, 'neigh_op_tnr_7')
// (7, 9, 'neigh_op_rgt_7')
// (7, 10, 'neigh_op_bnr_7')
// (8, 8, 'local_g1_7')
// (8, 8, 'lutff_5/in_3')
// (8, 8, 'neigh_op_top_7')
// (8, 9, 'lutff_7/out')
// (8, 10, 'neigh_op_bot_7')
// (9, 8, 'neigh_op_tnl_7')
// (9, 9, 'neigh_op_lft_7')
// (9, 10, 'neigh_op_bnl_7')

reg n459 = 0;
// (7, 8, 'sp12_h_r_0')
// (8, 7, 'neigh_op_tnr_6')
// (8, 8, 'neigh_op_rgt_6')
// (8, 8, 'sp12_h_r_3')
// (8, 9, 'neigh_op_bnr_6')
// (9, 7, 'neigh_op_top_6')
// (9, 8, 'lutff_6/out')
// (9, 8, 'sp12_h_r_4')
// (9, 9, 'neigh_op_bot_6')
// (10, 7, 'neigh_op_tnl_6')
// (10, 8, 'neigh_op_lft_6')
// (10, 8, 'sp12_h_r_7')
// (10, 9, 'neigh_op_bnl_6')
// (11, 8, 'local_g1_0')
// (11, 8, 'lutff_1/in_0')
// (11, 8, 'sp12_h_r_8')
// (12, 8, 'sp12_h_r_11')
// (13, 8, 'span12_horz_11')

reg n460 = 0;
// (7, 8, 'sp4_r_v_b_42')
// (7, 9, 'local_g1_7')
// (7, 9, 'lutff_0/in_2')
// (7, 9, 'lutff_6/in_2')
// (7, 9, 'sp4_r_v_b_31')
// (7, 10, 'sp4_r_v_b_18')
// (7, 11, 'sp4_r_v_b_7')
// (8, 6, 'neigh_op_tnr_6')
// (8, 7, 'neigh_op_rgt_6')
// (8, 7, 'sp4_h_r_1')
// (8, 7, 'sp4_v_t_42')
// (8, 8, 'neigh_op_bnr_6')
// (8, 8, 'sp4_v_b_42')
// (8, 9, 'sp4_v_b_31')
// (8, 10, 'sp4_v_b_18')
// (8, 11, 'sp4_v_b_7')
// (9, 6, 'neigh_op_top_6')
// (9, 7, 'lutff_6/out')
// (9, 7, 'sp4_h_r_12')
// (9, 7, 'sp4_r_v_b_45')
// (9, 8, 'neigh_op_bot_6')
// (9, 8, 'sp4_r_v_b_32')
// (9, 9, 'sp4_r_v_b_21')
// (9, 10, 'sp4_r_v_b_8')
// (10, 6, 'neigh_op_tnl_6')
// (10, 6, 'sp4_v_t_45')
// (10, 7, 'neigh_op_lft_6')
// (10, 7, 'sp4_h_r_25')
// (10, 7, 'sp4_v_b_45')
// (10, 8, 'neigh_op_bnl_6')
// (10, 8, 'sp4_v_b_32')
// (10, 9, 'sp4_v_b_21')
// (10, 10, 'sp4_h_r_8')
// (10, 10, 'sp4_v_b_8')
// (11, 4, 'sp4_r_v_b_42')
// (11, 5, 'sp4_r_v_b_31')
// (11, 6, 'local_g3_2')
// (11, 6, 'lutff_3/in_0')
// (11, 6, 'sp4_r_v_b_18')
// (11, 7, 'sp4_h_r_36')
// (11, 7, 'sp4_r_v_b_7')
// (11, 10, 'local_g0_5')
// (11, 10, 'lutff_3/in_0')
// (11, 10, 'sp4_h_r_21')
// (12, 3, 'sp4_v_t_42')
// (12, 4, 'sp4_v_b_42')
// (12, 5, 'sp4_v_b_31')
// (12, 6, 'sp4_v_b_18')
// (12, 7, 'sp4_h_l_36')
// (12, 7, 'sp4_v_b_7')
// (12, 10, 'sp4_h_r_32')
// (13, 10, 'span4_horz_32')

reg n461 = 0;
// (7, 8, 'sp4_r_v_b_43')
// (7, 9, 'local_g1_6')
// (7, 9, 'lutff_7/in_0')
// (7, 9, 'sp4_r_v_b_30')
// (7, 10, 'neigh_op_tnr_6')
// (7, 10, 'sp4_r_v_b_19')
// (7, 11, 'neigh_op_rgt_6')
// (7, 11, 'sp4_r_v_b_6')
// (7, 12, 'neigh_op_bnr_6')
// (8, 5, 'sp12_v_t_23')
// (8, 6, 'sp12_v_b_23')
// (8, 7, 'sp12_v_b_20')
// (8, 7, 'sp4_v_t_43')
// (8, 8, 'sp12_v_b_19')
// (8, 8, 'sp4_v_b_43')
// (8, 9, 'local_g2_0')
// (8, 9, 'local_g3_0')
// (8, 9, 'lutff_0/in_0')
// (8, 9, 'lutff_3/in_0')
// (8, 9, 'sp12_v_b_16')
// (8, 9, 'sp4_v_b_30')
// (8, 10, 'neigh_op_top_6')
// (8, 10, 'sp12_v_b_15')
// (8, 10, 'sp4_v_b_19')
// (8, 11, 'local_g1_6')
// (8, 11, 'lutff_6/out')
// (8, 11, 'lutff_7/in_0')
// (8, 11, 'sp12_v_b_12')
// (8, 11, 'sp4_v_b_6')
// (8, 12, 'neigh_op_bot_6')
// (8, 12, 'sp12_v_b_11')
// (8, 13, 'sp12_v_b_8')
// (8, 14, 'sp12_v_b_7')
// (8, 15, 'sp12_v_b_4')
// (8, 16, 'sp12_v_b_3')
// (8, 17, 'span12_vert_0')
// (9, 10, 'neigh_op_tnl_6')
// (9, 11, 'neigh_op_lft_6')
// (9, 12, 'neigh_op_bnl_6')

reg n462 = 0;
// (7, 9, 'neigh_op_tnr_0')
// (7, 10, 'neigh_op_rgt_0')
// (7, 11, 'neigh_op_bnr_0')
// (8, 9, 'neigh_op_top_0')
// (8, 10, 'local_g0_0')
// (8, 10, 'lutff_0/out')
// (8, 10, 'lutff_2/in_0')
// (8, 11, 'neigh_op_bot_0')
// (9, 9, 'neigh_op_tnl_0')
// (9, 10, 'neigh_op_lft_0')
// (9, 11, 'neigh_op_bnl_0')

reg n463 = 0;
// (7, 9, 'neigh_op_tnr_1')
// (7, 9, 'sp4_r_v_b_47')
// (7, 10, 'neigh_op_rgt_1')
// (7, 10, 'sp4_r_v_b_34')
// (7, 11, 'neigh_op_bnr_1')
// (7, 11, 'sp4_r_v_b_23')
// (7, 12, 'sp4_r_v_b_10')
// (8, 8, 'sp4_v_t_47')
// (8, 9, 'local_g2_7')
// (8, 9, 'lutff_6/in_3')
// (8, 9, 'neigh_op_top_1')
// (8, 9, 'sp4_v_b_47')
// (8, 10, 'lutff_1/out')
// (8, 10, 'sp4_v_b_34')
// (8, 11, 'neigh_op_bot_1')
// (8, 11, 'sp4_v_b_23')
// (8, 12, 'sp4_v_b_10')
// (9, 9, 'neigh_op_tnl_1')
// (9, 10, 'neigh_op_lft_1')
// (9, 11, 'neigh_op_bnl_1')

reg n464 = 0;
// (7, 9, 'neigh_op_tnr_2')
// (7, 10, 'neigh_op_rgt_2')
// (7, 11, 'neigh_op_bnr_2')
// (8, 9, 'neigh_op_top_2')
// (8, 10, 'local_g1_2')
// (8, 10, 'lutff_2/out')
// (8, 10, 'lutff_5/in_0')
// (8, 11, 'neigh_op_bot_2')
// (9, 9, 'neigh_op_tnl_2')
// (9, 10, 'neigh_op_lft_2')
// (9, 11, 'neigh_op_bnl_2')

reg n465 = 0;
// (7, 9, 'neigh_op_tnr_3')
// (7, 10, 'neigh_op_rgt_3')
// (7, 11, 'neigh_op_bnr_3')
// (8, 9, 'neigh_op_top_3')
// (8, 10, 'local_g0_3')
// (8, 10, 'lutff_1/in_0')
// (8, 10, 'lutff_3/out')
// (8, 11, 'neigh_op_bot_3')
// (9, 9, 'neigh_op_tnl_3')
// (9, 10, 'neigh_op_lft_3')
// (9, 11, 'neigh_op_bnl_3')

reg n466 = 0;
// (7, 9, 'neigh_op_tnr_4')
// (7, 10, 'neigh_op_rgt_4')
// (7, 11, 'neigh_op_bnr_4')
// (8, 9, 'neigh_op_top_4')
// (8, 10, 'local_g0_4')
// (8, 10, 'lutff_0/in_0')
// (8, 10, 'lutff_4/out')
// (8, 11, 'neigh_op_bot_4')
// (9, 9, 'neigh_op_tnl_4')
// (9, 10, 'neigh_op_lft_4')
// (9, 11, 'neigh_op_bnl_4')

reg n467 = 0;
// (7, 9, 'neigh_op_tnr_5')
// (7, 10, 'neigh_op_rgt_5')
// (7, 11, 'neigh_op_bnr_5')
// (8, 9, 'local_g0_5')
// (8, 9, 'lutff_7/in_0')
// (8, 9, 'neigh_op_top_5')
// (8, 10, 'lutff_5/out')
// (8, 11, 'neigh_op_bot_5')
// (9, 9, 'neigh_op_tnl_5')
// (9, 10, 'neigh_op_lft_5')
// (9, 11, 'neigh_op_bnl_5')

reg n468 = 0;
// (7, 9, 'neigh_op_tnr_6')
// (7, 10, 'neigh_op_rgt_6')
// (7, 11, 'neigh_op_bnr_6')
// (8, 9, 'neigh_op_top_6')
// (8, 10, 'local_g0_6')
// (8, 10, 'lutff_4/in_0')
// (8, 10, 'lutff_6/out')
// (8, 11, 'neigh_op_bot_6')
// (9, 9, 'neigh_op_tnl_6')
// (9, 10, 'neigh_op_lft_6')
// (9, 11, 'neigh_op_bnl_6')

reg n469 = 0;
// (7, 10, 'neigh_op_tnr_0')
// (7, 11, 'neigh_op_rgt_0')
// (7, 12, 'neigh_op_bnr_0')
// (8, 10, 'neigh_op_top_0')
// (8, 11, 'local_g0_0')
// (8, 11, 'lutff_0/out')
// (8, 11, 'lutff_6/in_0')
// (8, 12, 'neigh_op_bot_0')
// (9, 10, 'neigh_op_tnl_0')
// (9, 11, 'neigh_op_lft_0')
// (9, 12, 'neigh_op_bnl_0')

reg n470 = 0;
// (7, 10, 'neigh_op_tnr_1')
// (7, 11, 'neigh_op_rgt_1')
// (7, 12, 'neigh_op_bnr_1')
// (8, 0, 'span12_vert_22')
// (8, 1, 'sp12_v_b_22')
// (8, 2, 'sp12_v_b_21')
// (8, 3, 'sp12_v_b_18')
// (8, 4, 'sp12_v_b_17')
// (8, 5, 'sp12_v_b_14')
// (8, 6, 'sp12_v_b_13')
// (8, 7, 'local_g3_2')
// (8, 7, 'lutff_0/in_3')
// (8, 7, 'sp12_v_b_10')
// (8, 8, 'sp12_v_b_9')
// (8, 9, 'sp12_v_b_6')
// (8, 10, 'neigh_op_top_1')
// (8, 10, 'sp12_v_b_5')
// (8, 11, 'lutff_1/out')
// (8, 11, 'sp12_v_b_2')
// (8, 12, 'neigh_op_bot_1')
// (8, 12, 'sp12_v_b_1')
// (9, 10, 'neigh_op_tnl_1')
// (9, 11, 'neigh_op_lft_1')
// (9, 12, 'neigh_op_bnl_1')

reg n471 = 0;
// (7, 10, 'neigh_op_tnr_3')
// (7, 11, 'neigh_op_rgt_3')
// (7, 12, 'neigh_op_bnr_3')
// (8, 10, 'neigh_op_top_3')
// (8, 11, 'local_g0_3')
// (8, 11, 'lutff_1/in_0')
// (8, 11, 'lutff_3/out')
// (8, 12, 'neigh_op_bot_3')
// (9, 10, 'neigh_op_tnl_3')
// (9, 11, 'neigh_op_lft_3')
// (9, 12, 'neigh_op_bnl_3')

reg n472 = 0;
// (7, 10, 'neigh_op_tnr_4')
// (7, 11, 'neigh_op_rgt_4')
// (7, 12, 'neigh_op_bnr_4')
// (8, 10, 'neigh_op_top_4')
// (8, 11, 'local_g2_4')
// (8, 11, 'lutff_0/in_0')
// (8, 11, 'lutff_4/out')
// (8, 12, 'neigh_op_bot_4')
// (9, 10, 'neigh_op_tnl_4')
// (9, 11, 'neigh_op_lft_4')
// (9, 12, 'neigh_op_bnl_4')

reg n473 = 0;
// (7, 10, 'neigh_op_tnr_7')
// (7, 11, 'neigh_op_rgt_7')
// (7, 12, 'neigh_op_bnr_7')
// (8, 10, 'neigh_op_top_7')
// (8, 11, 'local_g1_7')
// (8, 11, 'lutff_4/in_0')
// (8, 11, 'lutff_7/out')
// (8, 12, 'neigh_op_bot_7')
// (9, 10, 'neigh_op_tnl_7')
// (9, 11, 'neigh_op_lft_7')
// (9, 12, 'neigh_op_bnl_7')

reg n474 = 0;
// (7, 10, 'sp4_r_v_b_36')
// (7, 11, 'sp4_r_v_b_25')
// (7, 12, 'sp4_r_v_b_12')
// (7, 13, 'sp4_r_v_b_1')
// (8, 9, 'local_g0_7')
// (8, 9, 'lutff_1/in_0')
// (8, 9, 'sp4_h_r_7')
// (8, 9, 'sp4_v_t_36')
// (8, 10, 'sp4_v_b_36')
// (8, 11, 'local_g3_1')
// (8, 11, 'lutff_7/in_1')
// (8, 11, 'sp4_v_b_25')
// (8, 12, 'sp4_v_b_12')
// (8, 13, 'sp4_v_b_1')
// (9, 9, 'sp4_h_r_18')
// (10, 8, 'neigh_op_tnr_5')
// (10, 9, 'neigh_op_rgt_5')
// (10, 9, 'sp4_h_r_31')
// (10, 10, 'neigh_op_bnr_5')
// (11, 8, 'neigh_op_top_5')
// (11, 9, 'lutff_5/out')
// (11, 9, 'sp4_h_r_42')
// (11, 10, 'neigh_op_bot_5')
// (12, 8, 'neigh_op_tnl_5')
// (12, 9, 'neigh_op_lft_5')
// (12, 9, 'sp4_h_l_42')
// (12, 10, 'neigh_op_bnl_5')

reg n475 = 0;
// (7, 11, 'neigh_op_tnr_0')
// (7, 12, 'neigh_op_rgt_0')
// (7, 13, 'neigh_op_bnr_0')
// (8, 11, 'neigh_op_top_0')
// (8, 12, 'local_g0_0')
// (8, 12, 'lutff_0/out')
// (8, 12, 'lutff_2/in_0')
// (8, 13, 'neigh_op_bot_0')
// (9, 11, 'neigh_op_tnl_0')
// (9, 12, 'neigh_op_lft_0')
// (9, 13, 'neigh_op_bnl_0')

reg n476 = 0;
// (7, 11, 'neigh_op_tnr_1')
// (7, 12, 'neigh_op_rgt_1')
// (7, 13, 'neigh_op_bnr_1')
// (8, 11, 'neigh_op_top_1')
// (8, 12, 'local_g1_1')
// (8, 12, 'lutff_0/in_0')
// (8, 12, 'lutff_1/out')
// (8, 13, 'neigh_op_bot_1')
// (9, 11, 'neigh_op_tnl_1')
// (9, 12, 'neigh_op_lft_1')
// (9, 13, 'neigh_op_bnl_1')

reg n477 = 0;
// (7, 11, 'neigh_op_tnr_2')
// (7, 12, 'neigh_op_rgt_2')
// (7, 13, 'neigh_op_bnr_2')
// (8, 11, 'local_g1_2')
// (8, 11, 'lutff_3/in_0')
// (8, 11, 'neigh_op_top_2')
// (8, 12, 'lutff_2/out')
// (8, 13, 'neigh_op_bot_2')
// (9, 11, 'neigh_op_tnl_2')
// (9, 12, 'neigh_op_lft_2')
// (9, 13, 'neigh_op_bnl_2')

reg n478 = 0;
// (7, 11, 'neigh_op_tnr_4')
// (7, 12, 'neigh_op_rgt_4')
// (7, 13, 'neigh_op_bnr_4')
// (8, 11, 'neigh_op_top_4')
// (8, 12, 'local_g0_4')
// (8, 12, 'lutff_4/out')
// (8, 12, 'lutff_6/in_0')
// (8, 13, 'neigh_op_bot_4')
// (9, 11, 'neigh_op_tnl_4')
// (9, 12, 'neigh_op_lft_4')
// (9, 13, 'neigh_op_bnl_4')

reg n479 = 0;
// (7, 11, 'neigh_op_tnr_5')
// (7, 12, 'neigh_op_rgt_5')
// (7, 13, 'neigh_op_bnr_5')
// (8, 11, 'neigh_op_top_5')
// (8, 12, 'local_g0_5')
// (8, 12, 'lutff_1/in_0')
// (8, 12, 'lutff_5/out')
// (8, 13, 'neigh_op_bot_5')
// (9, 11, 'neigh_op_tnl_5')
// (9, 12, 'neigh_op_lft_5')
// (9, 13, 'neigh_op_bnl_5')

reg n480 = 0;
// (7, 11, 'neigh_op_tnr_6')
// (7, 12, 'neigh_op_rgt_6')
// (7, 13, 'neigh_op_bnr_6')
// (8, 11, 'neigh_op_top_6')
// (8, 12, 'local_g1_6')
// (8, 12, 'lutff_5/in_0')
// (8, 12, 'lutff_6/out')
// (8, 13, 'neigh_op_bot_6')
// (9, 11, 'neigh_op_tnl_6')
// (9, 12, 'neigh_op_lft_6')
// (9, 13, 'neigh_op_bnl_6')

reg n481 = 0;
// (7, 12, 'neigh_op_tnr_0')
// (7, 13, 'neigh_op_rgt_0')
// (7, 14, 'neigh_op_bnr_0')
// (8, 12, 'neigh_op_top_0')
// (8, 13, 'local_g1_0')
// (8, 13, 'lutff_0/out')
// (8, 13, 'lutff_5/in_0')
// (8, 14, 'neigh_op_bot_0')
// (9, 12, 'neigh_op_tnl_0')
// (9, 13, 'neigh_op_lft_0')
// (9, 14, 'neigh_op_bnl_0')

reg n482 = 0;
// (7, 12, 'neigh_op_tnr_1')
// (7, 13, 'neigh_op_rgt_1')
// (7, 14, 'neigh_op_bnr_1')
// (8, 12, 'neigh_op_top_1')
// (8, 13, 'local_g1_1')
// (8, 13, 'lutff_0/in_0')
// (8, 13, 'lutff_1/out')
// (8, 14, 'neigh_op_bot_1')
// (9, 12, 'neigh_op_tnl_1')
// (9, 13, 'neigh_op_lft_1')
// (9, 14, 'neigh_op_bnl_1')

reg n483 = 0;
// (7, 12, 'neigh_op_tnr_7')
// (7, 13, 'neigh_op_rgt_7')
// (7, 14, 'neigh_op_bnr_7')
// (8, 12, 'neigh_op_top_7')
// (8, 13, 'local_g1_7')
// (8, 13, 'lutff_4/in_0')
// (8, 13, 'lutff_7/out')
// (8, 14, 'neigh_op_bot_7')
// (9, 12, 'neigh_op_tnl_7')
// (9, 13, 'neigh_op_lft_7')
// (9, 14, 'neigh_op_bnl_7')

wire n484;
// (8, 1, 'sp4_r_v_b_43')
// (8, 2, 'local_g0_6')
// (8, 2, 'local_g1_6')
// (8, 2, 'lutff_0/in_3')
// (8, 2, 'lutff_3/in_1')
// (8, 2, 'lutff_5/in_3')
// (8, 2, 'sp4_r_v_b_30')
// (8, 3, 'neigh_op_tnr_3')
// (8, 3, 'sp4_r_v_b_19')
// (8, 4, 'neigh_op_rgt_3')
// (8, 4, 'sp4_r_v_b_6')
// (8, 5, 'neigh_op_bnr_3')
// (9, 0, 'span4_vert_43')
// (9, 1, 'sp4_v_b_43')
// (9, 2, 'sp4_v_b_30')
// (9, 3, 'neigh_op_top_3')
// (9, 3, 'sp4_v_b_19')
// (9, 4, 'lutff_3/out')
// (9, 4, 'sp4_v_b_6')
// (9, 5, 'neigh_op_bot_3')
// (10, 3, 'neigh_op_tnl_3')
// (10, 4, 'neigh_op_lft_3')
// (10, 5, 'neigh_op_bnl_3')

wire n485;
// (8, 2, 'sp4_r_v_b_38')
// (8, 3, 'local_g0_3')
// (8, 3, 'lutff_1/in_2')
// (8, 3, 'lutff_2/in_1')
// (8, 3, 'neigh_op_tnr_7')
// (8, 3, 'sp4_r_v_b_27')
// (8, 4, 'local_g2_7')
// (8, 4, 'lutff_1/in_2')
// (8, 4, 'neigh_op_rgt_7')
// (8, 4, 'sp4_r_v_b_14')
// (8, 5, 'neigh_op_bnr_7')
// (8, 5, 'sp4_r_v_b_3')
// (9, 1, 'sp4_v_t_38')
// (9, 2, 'sp4_v_b_38')
// (9, 3, 'local_g1_7')
// (9, 3, 'lutff_7/in_3')
// (9, 3, 'neigh_op_top_7')
// (9, 3, 'sp4_v_b_27')
// (9, 4, 'lutff_7/out')
// (9, 4, 'sp4_v_b_14')
// (9, 5, 'neigh_op_bot_7')
// (9, 5, 'sp4_v_b_3')
// (10, 3, 'neigh_op_tnl_7')
// (10, 4, 'neigh_op_lft_7')
// (10, 5, 'neigh_op_bnl_7')

wire n486;
// (8, 3, 'neigh_op_tnr_0')
// (8, 4, 'local_g2_0')
// (8, 4, 'lutff_4/in_2')
// (8, 4, 'neigh_op_rgt_0')
// (8, 5, 'neigh_op_bnr_0')
// (9, 3, 'neigh_op_top_0')
// (9, 4, 'local_g1_0')
// (9, 4, 'local_g2_0')
// (9, 4, 'lutff_0/out')
// (9, 4, 'lutff_3/in_3')
// (9, 4, 'lutff_6/in_1')
// (9, 5, 'neigh_op_bot_0')
// (10, 3, 'neigh_op_tnl_0')
// (10, 4, 'neigh_op_lft_0')
// (10, 5, 'neigh_op_bnl_0')

wire n487;
// (8, 3, 'neigh_op_tnr_5')
// (8, 4, 'local_g2_5')
// (8, 4, 'lutff_2/in_1')
// (8, 4, 'lutff_5/in_2')
// (8, 4, 'neigh_op_rgt_5')
// (8, 5, 'neigh_op_bnr_5')
// (9, 3, 'neigh_op_top_5')
// (9, 4, 'local_g1_5')
// (9, 4, 'lutff_0/in_0')
// (9, 4, 'lutff_5/out')
// (9, 5, 'neigh_op_bot_5')
// (10, 3, 'neigh_op_tnl_5')
// (10, 4, 'neigh_op_lft_5')
// (10, 5, 'neigh_op_bnl_5')

wire n488;
// (8, 4, 'local_g2_3')
// (8, 4, 'local_g3_3')
// (8, 4, 'lutff_1/in_3')
// (8, 4, 'lutff_4/in_3')
// (8, 4, 'neigh_op_tnr_3')
// (8, 5, 'neigh_op_rgt_3')
// (8, 6, 'neigh_op_bnr_3')
// (9, 4, 'neigh_op_top_3')
// (9, 5, 'lutff_3/out')
// (9, 6, 'neigh_op_bot_3')
// (10, 4, 'neigh_op_tnl_3')
// (10, 5, 'neigh_op_lft_3')
// (10, 6, 'neigh_op_bnl_3')

reg n489 = 0;
// (8, 4, 'local_g3_5')
// (8, 4, 'lutff_7/in_3')
// (8, 4, 'sp4_r_v_b_45')
// (8, 5, 'sp4_r_v_b_32')
// (8, 6, 'neigh_op_tnr_4')
// (8, 6, 'sp4_r_v_b_21')
// (8, 7, 'neigh_op_rgt_4')
// (8, 7, 'sp4_r_v_b_8')
// (8, 8, 'neigh_op_bnr_4')
// (9, 3, 'sp4_v_t_45')
// (9, 4, 'sp4_v_b_45')
// (9, 5, 'sp4_v_b_32')
// (9, 6, 'neigh_op_top_4')
// (9, 6, 'sp4_v_b_21')
// (9, 7, 'lutff_4/out')
// (9, 7, 'sp4_v_b_8')
// (9, 8, 'neigh_op_bot_4')
// (10, 6, 'neigh_op_tnl_4')
// (10, 7, 'neigh_op_lft_4')
// (10, 8, 'neigh_op_bnl_4')

wire n490;
// (8, 4, 'neigh_op_tnr_1')
// (8, 5, 'neigh_op_rgt_1')
// (8, 6, 'neigh_op_bnr_1')
// (9, 4, 'neigh_op_top_1')
// (9, 5, 'local_g2_1')
// (9, 5, 'lutff_1/out')
// (9, 5, 'lutff_2/in_3')
// (9, 6, 'neigh_op_bot_1')
// (10, 4, 'neigh_op_tnl_1')
// (10, 5, 'neigh_op_lft_1')
// (10, 6, 'neigh_op_bnl_1')

wire n491;
// (8, 4, 'neigh_op_tnr_4')
// (8, 5, 'neigh_op_rgt_4')
// (8, 6, 'neigh_op_bnr_4')
// (9, 4, 'local_g0_4')
// (9, 4, 'lutff_3/in_1')
// (9, 4, 'neigh_op_top_4')
// (9, 5, 'local_g0_4')
// (9, 5, 'lutff_3/in_1')
// (9, 5, 'lutff_4/out')
// (9, 6, 'neigh_op_bot_4')
// (10, 4, 'neigh_op_tnl_4')
// (10, 5, 'neigh_op_lft_4')
// (10, 6, 'neigh_op_bnl_4')

wire n492;
// (8, 4, 'neigh_op_tnr_5')
// (8, 5, 'neigh_op_rgt_5')
// (8, 6, 'neigh_op_bnr_5')
// (9, 4, 'neigh_op_top_5')
// (9, 5, 'local_g0_5')
// (9, 5, 'local_g1_5')
// (9, 5, 'lutff_3/in_0')
// (9, 5, 'lutff_5/out')
// (9, 5, 'lutff_6/in_2')
// (9, 6, 'neigh_op_bot_5')
// (10, 4, 'neigh_op_tnl_5')
// (10, 5, 'neigh_op_lft_5')
// (10, 6, 'neigh_op_bnl_5')

wire n493;
// (8, 4, 'neigh_op_tnr_6')
// (8, 5, 'neigh_op_rgt_6')
// (8, 6, 'neigh_op_bnr_6')
// (9, 4, 'local_g1_6')
// (9, 4, 'lutff_6/in_3')
// (9, 4, 'neigh_op_top_6')
// (9, 5, 'lutff_6/out')
// (9, 6, 'neigh_op_bot_6')
// (10, 4, 'neigh_op_tnl_6')
// (10, 5, 'neigh_op_lft_6')
// (10, 6, 'neigh_op_bnl_6')

reg n494 = 0;
// (8, 4, 'neigh_op_tnr_7')
// (8, 5, 'neigh_op_rgt_7')
// (8, 6, 'neigh_op_bnr_7')
// (9, 4, 'neigh_op_top_7')
// (9, 5, 'local_g2_7')
// (9, 5, 'lutff_2/in_1')
// (9, 5, 'lutff_7/out')
// (9, 6, 'neigh_op_bot_7')
// (10, 4, 'neigh_op_tnl_7')
// (10, 5, 'neigh_op_lft_7')
// (10, 6, 'neigh_op_bnl_7')

wire n495;
// (8, 4, 'sp4_h_r_9')
// (9, 4, 'local_g1_4')
// (9, 4, 'lutff_0/in_1')
// (9, 4, 'lutff_7/in_2')
// (9, 4, 'sp4_h_r_20')
// (10, 3, 'neigh_op_tnr_6')
// (10, 4, 'neigh_op_rgt_6')
// (10, 4, 'sp4_h_r_33')
// (10, 5, 'neigh_op_bnr_6')
// (11, 3, 'neigh_op_top_6')
// (11, 4, 'lutff_6/out')
// (11, 4, 'sp4_h_r_44')
// (11, 5, 'neigh_op_bot_6')
// (12, 3, 'neigh_op_tnl_6')
// (12, 4, 'neigh_op_lft_6')
// (12, 4, 'sp4_h_l_44')
// (12, 5, 'neigh_op_bnl_6')

reg n496 = 0;
// (8, 4, 'sp4_r_v_b_38')
// (8, 5, 'sp4_r_v_b_27')
// (8, 6, 'sp4_r_v_b_14')
// (8, 7, 'sp4_r_v_b_3')
// (9, 3, 'sp4_v_t_38')
// (9, 4, 'sp4_v_b_38')
// (9, 5, 'local_g2_3')
// (9, 5, 'lutff_4/in_3')
// (9, 5, 'sp4_v_b_27')
// (9, 6, 'sp4_v_b_14')
// (9, 7, 'local_g0_2')
// (9, 7, 'lutff_6/in_0')
// (9, 7, 'sp4_h_r_10')
// (9, 7, 'sp4_v_b_3')
// (10, 6, 'neigh_op_tnr_1')
// (10, 7, 'neigh_op_rgt_1')
// (10, 7, 'sp4_h_r_23')
// (10, 8, 'neigh_op_bnr_1')
// (11, 6, 'neigh_op_top_1')
// (11, 7, 'lutff_1/out')
// (11, 7, 'sp4_h_r_34')
// (11, 8, 'neigh_op_bot_1')
// (12, 6, 'neigh_op_tnl_1')
// (12, 7, 'neigh_op_lft_1')
// (12, 7, 'sp4_h_r_47')
// (12, 8, 'neigh_op_bnl_1')
// (13, 7, 'span4_horz_47')

reg n497 = 0;
// (8, 4, 'sp4_r_v_b_39')
// (8, 5, 'sp4_r_v_b_26')
// (8, 6, 'sp4_r_v_b_15')
// (8, 7, 'local_g1_2')
// (8, 7, 'lutff_5/in_0')
// (8, 7, 'sp4_r_v_b_2')
// (8, 8, 'neigh_op_tnr_7')
// (8, 8, 'sp4_r_v_b_43')
// (8, 9, 'neigh_op_rgt_7')
// (8, 9, 'sp4_r_v_b_30')
// (8, 10, 'neigh_op_bnr_7')
// (8, 10, 'sp4_r_v_b_19')
// (8, 11, 'sp4_r_v_b_6')
// (9, 3, 'sp4_v_t_39')
// (9, 4, 'sp4_v_b_39')
// (9, 5, 'sp4_v_b_26')
// (9, 6, 'sp4_v_b_15')
// (9, 7, 'sp4_v_b_2')
// (9, 7, 'sp4_v_t_43')
// (9, 8, 'neigh_op_top_7')
// (9, 8, 'sp4_v_b_43')
// (9, 9, 'lutff_7/out')
// (9, 9, 'sp4_v_b_30')
// (9, 10, 'neigh_op_bot_7')
// (9, 10, 'sp4_v_b_19')
// (9, 11, 'sp4_v_b_6')
// (10, 8, 'neigh_op_tnl_7')
// (10, 9, 'neigh_op_lft_7')
// (10, 10, 'neigh_op_bnl_7')

reg n498 = 0;
// (8, 4, 'sp4_r_v_b_40')
// (8, 5, 'sp4_r_v_b_29')
// (8, 6, 'sp4_r_v_b_16')
// (8, 7, 'sp4_r_v_b_5')
// (8, 8, 'sp4_r_v_b_39')
// (8, 9, 'sp4_r_v_b_26')
// (8, 10, 'neigh_op_tnr_1')
// (8, 10, 'sp4_r_v_b_15')
// (8, 11, 'neigh_op_rgt_1')
// (8, 11, 'sp4_r_v_b_2')
// (8, 12, 'neigh_op_bnr_1')
// (9, 3, 'sp4_v_t_40')
// (9, 4, 'sp4_v_b_40')
// (9, 5, 'sp4_v_b_29')
// (9, 6, 'sp4_v_b_16')
// (9, 7, 'local_g0_5')
// (9, 7, 'lutff_0/in_3')
// (9, 7, 'sp4_v_b_5')
// (9, 7, 'sp4_v_t_39')
// (9, 8, 'sp4_v_b_39')
// (9, 9, 'sp4_v_b_26')
// (9, 10, 'neigh_op_top_1')
// (9, 10, 'sp4_v_b_15')
// (9, 11, 'lutff_1/out')
// (9, 11, 'sp4_v_b_2')
// (9, 12, 'neigh_op_bot_1')
// (10, 10, 'neigh_op_tnl_1')
// (10, 11, 'neigh_op_lft_1')
// (10, 12, 'neigh_op_bnl_1')

wire n499;
// (8, 5, 'local_g0_1')
// (8, 5, 'lutff_3/in_2')
// (8, 5, 'sp4_h_r_1')
// (9, 5, 'sp4_h_r_12')
// (10, 4, 'neigh_op_tnr_0')
// (10, 5, 'neigh_op_rgt_0')
// (10, 5, 'sp4_h_r_25')
// (10, 6, 'neigh_op_bnr_0')
// (11, 2, 'sp4_r_v_b_36')
// (11, 3, 'sp4_r_v_b_25')
// (11, 4, 'neigh_op_top_0')
// (11, 4, 'sp4_r_v_b_12')
// (11, 5, 'lutff_0/out')
// (11, 5, 'sp4_h_r_36')
// (11, 5, 'sp4_r_v_b_1')
// (11, 6, 'neigh_op_bot_0')
// (12, 1, 'sp4_v_t_36')
// (12, 2, 'sp4_v_b_36')
// (12, 3, 'sp4_v_b_25')
// (12, 4, 'neigh_op_tnl_0')
// (12, 4, 'sp4_v_b_12')
// (12, 5, 'neigh_op_lft_0')
// (12, 5, 'sp4_h_l_36')
// (12, 5, 'sp4_v_b_1')
// (12, 6, 'neigh_op_bnl_0')

reg n500 = 0;
// (8, 5, 'neigh_op_tnr_0')
// (8, 6, 'neigh_op_rgt_0')
// (8, 7, 'neigh_op_bnr_0')
// (9, 3, 'sp4_r_v_b_36')
// (9, 4, 'local_g1_1')
// (9, 4, 'lutff_5/in_3')
// (9, 4, 'sp4_r_v_b_25')
// (9, 5, 'neigh_op_top_0')
// (9, 5, 'sp4_r_v_b_12')
// (9, 6, 'local_g0_0')
// (9, 6, 'lutff_0/out')
// (9, 6, 'lutff_2/in_0')
// (9, 6, 'sp4_r_v_b_1')
// (9, 7, 'neigh_op_bot_0')
// (10, 2, 'sp4_v_t_36')
// (10, 3, 'sp4_v_b_36')
// (10, 4, 'sp4_v_b_25')
// (10, 5, 'neigh_op_tnl_0')
// (10, 5, 'sp4_v_b_12')
// (10, 6, 'neigh_op_lft_0')
// (10, 6, 'sp4_v_b_1')
// (10, 7, 'neigh_op_bnl_0')

reg n501 = 0;
// (8, 5, 'neigh_op_tnr_4')
// (8, 6, 'neigh_op_rgt_4')
// (8, 7, 'neigh_op_bnr_4')
// (9, 5, 'neigh_op_top_4')
// (9, 6, 'local_g0_4')
// (9, 6, 'lutff_0/in_0')
// (9, 6, 'lutff_4/out')
// (9, 7, 'neigh_op_bot_4')
// (10, 5, 'neigh_op_tnl_4')
// (10, 6, 'neigh_op_lft_4')
// (10, 7, 'neigh_op_bnl_4')

reg n502 = 0;
// (8, 5, 'neigh_op_tnr_5')
// (8, 6, 'neigh_op_rgt_5')
// (8, 7, 'neigh_op_bnr_5')
// (9, 5, 'neigh_op_top_5')
// (9, 6, 'local_g2_5')
// (9, 6, 'lutff_1/in_0')
// (9, 6, 'lutff_5/out')
// (9, 7, 'neigh_op_bot_5')
// (10, 5, 'neigh_op_tnl_5')
// (10, 6, 'neigh_op_lft_5')
// (10, 7, 'neigh_op_bnl_5')

reg n503 = 0;
// (8, 5, 'neigh_op_tnr_7')
// (8, 6, 'neigh_op_rgt_7')
// (8, 7, 'neigh_op_bnr_7')
// (9, 5, 'neigh_op_top_7')
// (9, 6, 'local_g1_7')
// (9, 6, 'lutff_5/in_3')
// (9, 6, 'lutff_7/out')
// (9, 7, 'neigh_op_bot_7')
// (10, 5, 'neigh_op_tnl_7')
// (10, 6, 'neigh_op_lft_7')
// (10, 7, 'neigh_op_bnl_7')

reg n504 = 0;
// (8, 6, 'neigh_op_tnr_0')
// (8, 7, 'neigh_op_rgt_0')
// (8, 8, 'neigh_op_bnr_0')
// (9, 6, 'neigh_op_top_0')
// (9, 7, 'local_g1_0')
// (9, 7, 'lutff_0/out')
// (9, 7, 'lutff_5/in_0')
// (9, 8, 'neigh_op_bot_0')
// (10, 6, 'neigh_op_tnl_0')
// (10, 7, 'neigh_op_lft_0')
// (10, 8, 'neigh_op_bnl_0')

reg n505 = 0;
// (8, 6, 'neigh_op_tnr_2')
// (8, 7, 'neigh_op_rgt_2')
// (8, 8, 'neigh_op_bnr_2')
// (9, 6, 'neigh_op_top_2')
// (9, 7, 'local_g1_2')
// (9, 7, 'lutff_2/out')
// (9, 7, 'lutff_7/in_0')
// (9, 8, 'neigh_op_bot_2')
// (10, 6, 'neigh_op_tnl_2')
// (10, 7, 'neigh_op_lft_2')
// (10, 8, 'neigh_op_bnl_2')

reg n506 = 0;
// (8, 6, 'neigh_op_tnr_5')
// (8, 7, 'local_g2_5')
// (8, 7, 'lutff_7/in_0')
// (8, 7, 'neigh_op_rgt_5')
// (8, 8, 'neigh_op_bnr_5')
// (9, 6, 'neigh_op_top_5')
// (9, 7, 'lutff_5/out')
// (9, 8, 'neigh_op_bot_5')
// (10, 6, 'neigh_op_tnl_5')
// (10, 7, 'neigh_op_lft_5')
// (10, 8, 'neigh_op_bnl_5')

reg n507 = 0;
// (8, 6, 'neigh_op_tnr_7')
// (8, 7, 'neigh_op_rgt_7')
// (8, 8, 'neigh_op_bnr_7')
// (9, 2, 'sp12_v_t_22')
// (9, 3, 'sp12_v_b_22')
// (9, 4, 'sp12_v_b_21')
// (9, 5, 'local_g2_2')
// (9, 5, 'lutff_2/in_2')
// (9, 5, 'sp12_v_b_18')
// (9, 6, 'neigh_op_top_7')
// (9, 6, 'sp12_v_b_17')
// (9, 7, 'local_g0_7')
// (9, 7, 'lutff_3/in_0')
// (9, 7, 'lutff_7/out')
// (9, 7, 'sp12_v_b_14')
// (9, 8, 'neigh_op_bot_7')
// (9, 8, 'sp12_v_b_13')
// (9, 9, 'sp12_v_b_10')
// (9, 10, 'sp12_v_b_9')
// (9, 11, 'sp12_v_b_6')
// (9, 12, 'sp12_v_b_5')
// (9, 13, 'sp12_v_b_2')
// (9, 14, 'sp12_v_b_1')
// (10, 6, 'neigh_op_tnl_7')
// (10, 7, 'neigh_op_lft_7')
// (10, 8, 'neigh_op_bnl_7')

wire \d_out[3] ;
// (8, 7, 'neigh_op_tnr_1')
// (8, 8, 'neigh_op_rgt_1')
// (8, 8, 'sp4_h_r_7')
// (8, 9, 'neigh_op_bnr_1')
// (9, 7, 'neigh_op_top_1')
// (9, 8, 'lutff_1/out')
// (9, 8, 'sp4_h_r_18')
// (9, 9, 'neigh_op_bot_1')
// (10, 7, 'neigh_op_tnl_1')
// (10, 8, 'neigh_op_lft_1')
// (10, 8, 'sp4_h_r_31')
// (10, 9, 'neigh_op_bnl_1')
// (11, 8, 'sp4_h_r_42')
// (12, 8, 'sp4_h_l_42')
// (12, 8, 'sp4_h_r_7')
// (13, 8, 'span4_horz_7')
// (13, 8, 'span4_vert_t_13')
// (13, 9, 'span4_vert_b_13')
// (13, 10, 'span4_vert_b_9')
// (13, 11, 'io_0/D_OUT_0')
// (13, 11, 'io_0/PAD')
// (13, 11, 'local_g1_5')
// (13, 11, 'span4_vert_b_5')
// (13, 12, 'span4_vert_b_1')

reg n509 = 0;
// (8, 7, 'neigh_op_tnr_3')
// (8, 8, 'neigh_op_rgt_3')
// (8, 9, 'neigh_op_bnr_3')
// (9, 0, 'span12_vert_21')
// (9, 1, 'sp12_v_b_21')
// (9, 2, 'sp12_v_b_18')
// (9, 3, 'sp12_v_b_17')
// (9, 4, 'sp12_v_b_14')
// (9, 5, 'sp12_v_b_13')
// (9, 6, 'local_g2_2')
// (9, 6, 'lutff_4/in_0')
// (9, 6, 'sp12_v_b_10')
// (9, 7, 'neigh_op_top_3')
// (9, 7, 'sp12_v_b_9')
// (9, 8, 'lutff_3/out')
// (9, 8, 'sp12_v_b_6')
// (9, 9, 'neigh_op_bot_3')
// (9, 9, 'sp12_v_b_5')
// (9, 10, 'sp12_v_b_2')
// (9, 11, 'sp12_v_b_1')
// (10, 7, 'neigh_op_tnl_3')
// (10, 8, 'neigh_op_lft_3')
// (10, 9, 'neigh_op_bnl_3')

reg n510 = 0;
// (8, 7, 'neigh_op_tnr_5')
// (8, 8, 'neigh_op_rgt_5')
// (8, 9, 'neigh_op_bnr_5')
// (9, 7, 'local_g1_5')
// (9, 7, 'lutff_2/in_0')
// (9, 7, 'neigh_op_top_5')
// (9, 8, 'lutff_5/out')
// (9, 9, 'neigh_op_bot_5')
// (10, 7, 'neigh_op_tnl_5')
// (10, 8, 'neigh_op_lft_5')
// (10, 9, 'neigh_op_bnl_5')

reg n511 = 0;
// (8, 7, 'sp4_h_r_2')
// (9, 7, 'local_g1_7')
// (9, 7, 'lutff_4/in_0')
// (9, 7, 'sp4_h_r_15')
// (10, 7, 'neigh_op_tnr_3')
// (10, 7, 'sp4_h_r_26')
// (10, 8, 'neigh_op_rgt_3')
// (10, 9, 'neigh_op_bnr_3')
// (11, 7, 'neigh_op_top_3')
// (11, 7, 'sp4_h_r_39')
// (11, 8, 'lutff_3/out')
// (11, 8, 'sp4_r_v_b_39')
// (11, 9, 'neigh_op_bot_3')
// (11, 9, 'sp4_r_v_b_26')
// (11, 10, 'sp4_r_v_b_15')
// (11, 11, 'sp4_r_v_b_2')
// (12, 7, 'neigh_op_tnl_3')
// (12, 7, 'sp4_h_l_39')
// (12, 7, 'sp4_v_t_39')
// (12, 8, 'neigh_op_lft_3')
// (12, 8, 'sp4_v_b_39')
// (12, 9, 'neigh_op_bnl_3')
// (12, 9, 'sp4_v_b_26')
// (12, 10, 'sp4_v_b_15')
// (12, 11, 'sp4_v_b_2')

reg n512 = 0;
// (8, 8, 'neigh_op_tnr_0')
// (8, 9, 'neigh_op_rgt_0')
// (8, 10, 'neigh_op_bnr_0')
// (9, 0, 'span12_vert_16')
// (9, 1, 'sp12_v_b_16')
// (9, 2, 'sp12_v_b_15')
// (9, 3, 'sp12_v_b_12')
// (9, 4, 'sp12_v_b_11')
// (9, 5, 'sp12_v_b_8')
// (9, 6, 'local_g2_7')
// (9, 6, 'lutff_7/in_0')
// (9, 6, 'sp12_v_b_7')
// (9, 7, 'sp12_v_b_4')
// (9, 8, 'neigh_op_top_0')
// (9, 8, 'sp12_v_b_3')
// (9, 9, 'lutff_0/out')
// (9, 9, 'sp12_v_b_0')
// (9, 10, 'neigh_op_bot_0')
// (10, 8, 'neigh_op_tnl_0')
// (10, 9, 'neigh_op_lft_0')
// (10, 10, 'neigh_op_bnl_0')

reg n513 = 0;
// (8, 8, 'neigh_op_tnr_2')
// (8, 9, 'neigh_op_rgt_2')
// (8, 10, 'neigh_op_bnr_2')
// (9, 8, 'neigh_op_top_2')
// (9, 9, 'local_g0_2')
// (9, 9, 'lutff_2/out')
// (9, 9, 'lutff_5/in_3')
// (9, 10, 'neigh_op_bot_2')
// (10, 8, 'neigh_op_tnl_2')
// (10, 9, 'neigh_op_lft_2')
// (10, 10, 'neigh_op_bnl_2')

reg n514 = 0;
// (8, 8, 'neigh_op_tnr_3')
// (8, 9, 'neigh_op_rgt_3')
// (8, 10, 'neigh_op_bnr_3')
// (9, 8, 'neigh_op_top_3')
// (9, 9, 'local_g3_3')
// (9, 9, 'lutff_0/in_0')
// (9, 9, 'lutff_3/out')
// (9, 10, 'neigh_op_bot_3')
// (10, 8, 'neigh_op_tnl_3')
// (10, 9, 'neigh_op_lft_3')
// (10, 10, 'neigh_op_bnl_3')

reg n515 = 0;
// (8, 8, 'neigh_op_tnr_5')
// (8, 9, 'neigh_op_rgt_5')
// (8, 10, 'neigh_op_bnr_5')
// (9, 8, 'neigh_op_top_5')
// (9, 9, 'local_g0_5')
// (9, 9, 'lutff_5/out')
// (9, 9, 'lutff_7/in_0')
// (9, 10, 'neigh_op_bot_5')
// (10, 8, 'neigh_op_tnl_5')
// (10, 9, 'neigh_op_lft_5')
// (10, 10, 'neigh_op_bnl_5')

reg n516 = 0;
// (8, 8, 'neigh_op_tnr_6')
// (8, 9, 'neigh_op_rgt_6')
// (8, 10, 'neigh_op_bnr_6')
// (9, 8, 'neigh_op_top_6')
// (9, 9, 'local_g1_6')
// (9, 9, 'lutff_1/in_0')
// (9, 9, 'lutff_6/out')
// (9, 10, 'neigh_op_bot_6')
// (10, 8, 'neigh_op_tnl_6')
// (10, 9, 'neigh_op_lft_6')
// (10, 10, 'neigh_op_bnl_6')

reg n517 = 0;
// (8, 9, 'neigh_op_tnr_1')
// (8, 10, 'neigh_op_rgt_1')
// (8, 11, 'neigh_op_bnr_1')
// (9, 9, 'neigh_op_top_1')
// (9, 10, 'local_g0_1')
// (9, 10, 'lutff_1/out')
// (9, 10, 'lutff_5/in_0')
// (9, 11, 'neigh_op_bot_1')
// (10, 9, 'neigh_op_tnl_1')
// (10, 10, 'neigh_op_lft_1')
// (10, 11, 'neigh_op_bnl_1')

reg n518 = 0;
// (8, 9, 'neigh_op_tnr_2')
// (8, 10, 'neigh_op_rgt_2')
// (8, 11, 'neigh_op_bnr_2')
// (9, 9, 'neigh_op_top_2')
// (9, 10, 'local_g2_2')
// (9, 10, 'lutff_2/out')
// (9, 10, 'lutff_4/in_0')
// (9, 11, 'neigh_op_bot_2')
// (10, 9, 'neigh_op_tnl_2')
// (10, 10, 'neigh_op_lft_2')
// (10, 11, 'neigh_op_bnl_2')

reg n519 = 0;
// (8, 9, 'neigh_op_tnr_3')
// (8, 10, 'neigh_op_rgt_3')
// (8, 11, 'neigh_op_bnr_3')
// (9, 9, 'neigh_op_top_3')
// (9, 10, 'local_g0_3')
// (9, 10, 'lutff_1/in_0')
// (9, 10, 'lutff_3/out')
// (9, 11, 'neigh_op_bot_3')
// (10, 9, 'neigh_op_tnl_3')
// (10, 10, 'neigh_op_lft_3')
// (10, 11, 'neigh_op_bnl_3')

reg n520 = 0;
// (8, 9, 'neigh_op_tnr_4')
// (8, 10, 'neigh_op_rgt_4')
// (8, 11, 'neigh_op_bnr_4')
// (9, 9, 'local_g0_4')
// (9, 9, 'lutff_2/in_0')
// (9, 9, 'neigh_op_top_4')
// (9, 10, 'lutff_4/out')
// (9, 11, 'neigh_op_bot_4')
// (10, 9, 'neigh_op_tnl_4')
// (10, 10, 'neigh_op_lft_4')
// (10, 11, 'neigh_op_bnl_4')

reg n521 = 0;
// (8, 9, 'neigh_op_tnr_5')
// (8, 10, 'neigh_op_rgt_5')
// (8, 11, 'neigh_op_bnr_5')
// (9, 9, 'neigh_op_top_5')
// (9, 10, 'local_g1_5')
// (9, 10, 'lutff_2/in_0')
// (9, 10, 'lutff_5/out')
// (9, 11, 'neigh_op_bot_5')
// (10, 9, 'neigh_op_tnl_5')
// (10, 10, 'neigh_op_lft_5')
// (10, 11, 'neigh_op_bnl_5')

reg n522 = 0;
// (8, 9, 'neigh_op_tnr_7')
// (8, 10, 'neigh_op_rgt_7')
// (8, 10, 'sp4_h_r_3')
// (8, 11, 'neigh_op_bnr_7')
// (9, 9, 'neigh_op_top_7')
// (9, 10, 'lutff_7/out')
// (9, 10, 'sp4_h_r_14')
// (9, 11, 'neigh_op_bot_7')
// (10, 9, 'neigh_op_tnl_7')
// (10, 10, 'neigh_op_lft_7')
// (10, 10, 'sp4_h_r_27')
// (10, 11, 'neigh_op_bnl_7')
// (11, 10, 'local_g2_6')
// (11, 10, 'lutff_4/in_0')
// (11, 10, 'sp4_h_r_38')
// (12, 10, 'sp4_h_l_38')

reg n523 = 0;
// (8, 10, 'local_g1_1')
// (8, 10, 'lutff_6/in_0')
// (8, 10, 'sp4_h_r_9')
// (9, 10, 'sp4_h_r_20')
// (10, 9, 'neigh_op_tnr_6')
// (10, 10, 'neigh_op_rgt_6')
// (10, 10, 'sp4_h_r_33')
// (10, 11, 'neigh_op_bnr_6')
// (11, 9, 'neigh_op_top_6')
// (11, 10, 'lutff_6/out')
// (11, 10, 'sp4_h_r_44')
// (11, 11, 'neigh_op_bot_6')
// (12, 9, 'neigh_op_tnl_6')
// (12, 10, 'neigh_op_lft_6')
// (12, 10, 'sp4_h_l_44')
// (12, 11, 'neigh_op_bnl_6')

reg n524 = 0;
// (8, 10, 'neigh_op_tnr_2')
// (8, 11, 'neigh_op_rgt_2')
// (8, 12, 'neigh_op_bnr_2')
// (9, 1, 'sp12_v_t_23')
// (9, 2, 'sp12_v_b_23')
// (9, 3, 'sp12_v_b_20')
// (9, 4, 'sp12_v_b_19')
// (9, 5, 'local_g2_0')
// (9, 5, 'lutff_5/in_3')
// (9, 5, 'sp12_v_b_16')
// (9, 6, 'sp12_v_b_15')
// (9, 7, 'sp12_v_b_12')
// (9, 8, 'sp12_v_b_11')
// (9, 9, 'sp12_v_b_8')
// (9, 10, 'local_g0_2')
// (9, 10, 'lutff_0/in_0')
// (9, 10, 'neigh_op_top_2')
// (9, 10, 'sp12_v_b_7')
// (9, 11, 'lutff_2/out')
// (9, 11, 'sp12_v_b_4')
// (9, 12, 'neigh_op_bot_2')
// (9, 12, 'sp12_v_b_3')
// (9, 13, 'sp12_v_b_0')
// (10, 10, 'neigh_op_tnl_2')
// (10, 11, 'neigh_op_lft_2')
// (10, 12, 'neigh_op_bnl_2')

reg n525 = 0;
// (8, 10, 'neigh_op_tnr_5')
// (8, 11, 'neigh_op_rgt_5')
// (8, 12, 'neigh_op_bnr_5')
// (9, 10, 'neigh_op_top_5')
// (9, 11, 'local_g1_5')
// (9, 11, 'lutff_2/in_0')
// (9, 11, 'lutff_5/out')
// (9, 12, 'neigh_op_bot_5')
// (10, 10, 'neigh_op_tnl_5')
// (10, 11, 'neigh_op_lft_5')
// (10, 12, 'neigh_op_bnl_5')

reg n526 = 0;
// (8, 10, 'sp4_h_r_5')
// (9, 10, 'local_g1_0')
// (9, 10, 'lutff_3/in_0')
// (9, 10, 'sp4_h_r_16')
// (10, 9, 'neigh_op_tnr_4')
// (10, 10, 'neigh_op_rgt_4')
// (10, 10, 'sp4_h_r_29')
// (10, 11, 'neigh_op_bnr_4')
// (11, 9, 'neigh_op_top_4')
// (11, 10, 'lutff_4/out')
// (11, 10, 'sp4_h_r_40')
// (11, 11, 'neigh_op_bot_4')
// (12, 9, 'neigh_op_tnl_4')
// (12, 10, 'neigh_op_lft_4')
// (12, 10, 'sp4_h_l_40')
// (12, 11, 'neigh_op_bnl_4')

reg n527 = 0;
// (8, 11, 'neigh_op_tnr_0')
// (8, 12, 'neigh_op_rgt_0')
// (8, 13, 'neigh_op_bnr_0')
// (9, 11, 'neigh_op_top_0')
// (9, 12, 'local_g0_0')
// (9, 12, 'lutff_0/out')
// (9, 12, 'lutff_6/in_0')
// (9, 13, 'neigh_op_bot_0')
// (10, 11, 'neigh_op_tnl_0')
// (10, 12, 'neigh_op_lft_0')
// (10, 13, 'neigh_op_bnl_0')

reg n528 = 0;
// (8, 11, 'neigh_op_tnr_1')
// (8, 12, 'neigh_op_rgt_1')
// (8, 13, 'neigh_op_bnr_1')
// (9, 11, 'neigh_op_top_1')
// (9, 12, 'local_g0_1')
// (9, 12, 'lutff_1/out')
// (9, 12, 'lutff_3/in_0')
// (9, 13, 'neigh_op_bot_1')
// (10, 11, 'neigh_op_tnl_1')
// (10, 12, 'neigh_op_lft_1')
// (10, 13, 'neigh_op_bnl_1')

reg n529 = 0;
// (8, 11, 'neigh_op_tnr_3')
// (8, 12, 'neigh_op_rgt_3')
// (8, 12, 'sp4_h_r_11')
// (8, 13, 'neigh_op_bnr_3')
// (9, 11, 'neigh_op_top_3')
// (9, 12, 'lutff_3/out')
// (9, 12, 'sp4_h_r_22')
// (9, 13, 'neigh_op_bot_3')
// (10, 11, 'neigh_op_tnl_3')
// (10, 12, 'neigh_op_lft_3')
// (10, 12, 'sp4_h_r_35')
// (10, 13, 'neigh_op_bnl_3')
// (11, 12, 'local_g3_6')
// (11, 12, 'lutff_3/in_0')
// (11, 12, 'sp4_h_r_46')
// (12, 12, 'sp4_h_l_46')

reg n530 = 0;
// (8, 11, 'neigh_op_tnr_5')
// (8, 12, 'neigh_op_rgt_5')
// (8, 13, 'neigh_op_bnr_5')
// (9, 11, 'neigh_op_top_5')
// (9, 12, 'local_g0_5')
// (9, 12, 'lutff_1/in_0')
// (9, 12, 'lutff_5/out')
// (9, 13, 'neigh_op_bot_5')
// (10, 11, 'neigh_op_tnl_5')
// (10, 12, 'neigh_op_lft_5')
// (10, 13, 'neigh_op_bnl_5')

reg n531 = 0;
// (8, 11, 'neigh_op_tnr_6')
// (8, 12, 'neigh_op_rgt_6')
// (8, 13, 'neigh_op_bnr_6')
// (9, 11, 'local_g1_6')
// (9, 11, 'lutff_1/in_0')
// (9, 11, 'neigh_op_top_6')
// (9, 12, 'lutff_6/out')
// (9, 13, 'neigh_op_bot_6')
// (10, 11, 'neigh_op_tnl_6')
// (10, 12, 'neigh_op_lft_6')
// (10, 13, 'neigh_op_bnl_6')

reg n532 = 0;
// (8, 12, 'neigh_op_tnr_5')
// (8, 13, 'neigh_op_rgt_5')
// (8, 14, 'neigh_op_bnr_5')
// (9, 10, 'sp4_r_v_b_46')
// (9, 11, 'local_g2_3')
// (9, 11, 'lutff_5/in_0')
// (9, 11, 'sp4_r_v_b_35')
// (9, 12, 'neigh_op_top_5')
// (9, 12, 'sp4_r_v_b_22')
// (9, 13, 'lutff_5/out')
// (9, 13, 'sp4_r_v_b_11')
// (9, 14, 'neigh_op_bot_5')
// (10, 9, 'sp4_v_t_46')
// (10, 10, 'sp4_v_b_46')
// (10, 11, 'sp4_v_b_35')
// (10, 12, 'neigh_op_tnl_5')
// (10, 12, 'sp4_v_b_22')
// (10, 13, 'neigh_op_lft_5')
// (10, 13, 'sp4_v_b_11')
// (10, 14, 'neigh_op_bnl_5')

reg n533 = 0;
// (8, 12, 'sp4_h_r_1')
// (9, 12, 'local_g0_4')
// (9, 12, 'lutff_0/in_0')
// (9, 12, 'sp4_h_r_12')
// (10, 11, 'neigh_op_tnr_2')
// (10, 12, 'neigh_op_rgt_2')
// (10, 12, 'sp4_h_r_25')
// (10, 13, 'neigh_op_bnr_2')
// (11, 11, 'neigh_op_top_2')
// (11, 12, 'lutff_2/out')
// (11, 12, 'sp4_h_r_36')
// (11, 13, 'neigh_op_bot_2')
// (12, 11, 'neigh_op_tnl_2')
// (12, 12, 'neigh_op_lft_2')
// (12, 12, 'sp4_h_l_36')
// (12, 13, 'neigh_op_bnl_2')

reg n534 = 0;
// (10, 3, 'neigh_op_tnr_7')
// (10, 4, 'neigh_op_rgt_7')
// (10, 5, 'neigh_op_bnr_7')
// (11, 3, 'neigh_op_top_7')
// (11, 4, 'lutff_7/out')
// (11, 5, 'local_g0_7')
// (11, 5, 'lutff_7/in_0')
// (11, 5, 'neigh_op_bot_7')
// (12, 3, 'neigh_op_tnl_7')
// (12, 4, 'neigh_op_lft_7')
// (12, 5, 'neigh_op_bnl_7')

reg n535 = 0;
// (10, 4, 'neigh_op_tnr_7')
// (10, 5, 'neigh_op_rgt_7')
// (10, 6, 'neigh_op_bnr_7')
// (11, 4, 'neigh_op_top_7')
// (11, 5, 'local_g1_7')
// (11, 5, 'lutff_6/in_0')
// (11, 5, 'lutff_7/out')
// (11, 6, 'neigh_op_bot_7')
// (12, 4, 'neigh_op_tnl_7')
// (12, 5, 'neigh_op_lft_7')
// (12, 6, 'neigh_op_bnl_7')

reg n536 = 0;
// (10, 5, 'neigh_op_tnr_2')
// (10, 6, 'neigh_op_rgt_2')
// (10, 7, 'neigh_op_bnr_2')
// (11, 0, 'span12_vert_15')
// (11, 1, 'sp12_v_b_15')
// (11, 2, 'sp12_v_b_12')
// (11, 3, 'sp12_v_b_11')
// (11, 4, 'local_g3_0')
// (11, 4, 'lutff_2/in_3')
// (11, 4, 'sp12_v_b_8')
// (11, 5, 'neigh_op_top_2')
// (11, 5, 'sp12_v_b_7')
// (11, 6, 'lutff_2/out')
// (11, 6, 'sp12_v_b_4')
// (11, 7, 'neigh_op_bot_2')
// (11, 7, 'sp12_v_b_3')
// (11, 8, 'sp12_v_b_0')
// (12, 5, 'neigh_op_tnl_2')
// (12, 6, 'neigh_op_lft_2')
// (12, 7, 'neigh_op_bnl_2')

reg n537 = 0;
// (10, 5, 'neigh_op_tnr_3')
// (10, 6, 'neigh_op_rgt_3')
// (10, 7, 'neigh_op_bnr_3')
// (11, 5, 'local_g1_3')
// (11, 5, 'lutff_3/in_3')
// (11, 5, 'neigh_op_top_3')
// (11, 6, 'lutff_3/out')
// (11, 7, 'neigh_op_bot_3')
// (12, 5, 'neigh_op_tnl_3')
// (12, 6, 'neigh_op_lft_3')
// (12, 7, 'neigh_op_bnl_3')

reg n538 = 0;
// (10, 5, 'neigh_op_tnr_6')
// (10, 6, 'neigh_op_rgt_6')
// (10, 7, 'neigh_op_bnr_6')
// (11, 5, 'local_g0_6')
// (11, 5, 'lutff_1/in_3')
// (11, 5, 'neigh_op_top_6')
// (11, 6, 'lutff_6/out')
// (11, 7, 'neigh_op_bot_6')
// (12, 5, 'neigh_op_tnl_6')
// (12, 6, 'neigh_op_lft_6')
// (12, 7, 'neigh_op_bnl_6')

reg n539 = 0;
// (10, 6, 'neigh_op_tnr_0')
// (10, 7, 'neigh_op_rgt_0')
// (10, 8, 'neigh_op_bnr_0')
// (11, 6, 'neigh_op_top_0')
// (11, 7, 'lutff_0/out')
// (11, 8, 'neigh_op_bot_0')
// (12, 6, 'neigh_op_tnl_0')
// (12, 7, 'local_g0_0')
// (12, 7, 'lutff_2/in_0')
// (12, 7, 'neigh_op_lft_0')
// (12, 8, 'neigh_op_bnl_0')

reg n540 = 0;
// (10, 6, 'neigh_op_tnr_3')
// (10, 7, 'neigh_op_rgt_3')
// (10, 8, 'neigh_op_bnr_3')
// (11, 6, 'neigh_op_top_3')
// (11, 7, 'local_g1_3')
// (11, 7, 'lutff_3/out')
// (11, 7, 'lutff_4/in_0')
// (11, 8, 'neigh_op_bot_3')
// (12, 6, 'neigh_op_tnl_3')
// (12, 7, 'neigh_op_lft_3')
// (12, 8, 'neigh_op_bnl_3')

reg n541 = 0;
// (10, 6, 'neigh_op_tnr_4')
// (10, 7, 'neigh_op_rgt_4')
// (10, 8, 'neigh_op_bnr_4')
// (11, 6, 'neigh_op_top_4')
// (11, 7, 'local_g0_4')
// (11, 7, 'lutff_0/in_0')
// (11, 7, 'lutff_4/out')
// (11, 8, 'neigh_op_bot_4')
// (12, 6, 'neigh_op_tnl_4')
// (12, 7, 'neigh_op_lft_4')
// (12, 8, 'neigh_op_bnl_4')

reg n542 = 0;
// (10, 7, 'neigh_op_tnr_1')
// (10, 8, 'neigh_op_rgt_1')
// (10, 9, 'neigh_op_bnr_1')
// (11, 7, 'local_g0_1')
// (11, 7, 'lutff_1/in_0')
// (11, 7, 'neigh_op_top_1')
// (11, 8, 'lutff_1/out')
// (11, 9, 'neigh_op_bot_1')
// (12, 7, 'neigh_op_tnl_1')
// (12, 8, 'neigh_op_lft_1')
// (12, 9, 'neigh_op_bnl_1')

reg n543 = 0;
// (10, 8, 'neigh_op_tnr_3')
// (10, 9, 'neigh_op_rgt_3')
// (10, 10, 'neigh_op_bnr_3')
// (11, 8, 'neigh_op_top_3')
// (11, 9, 'lutff_3/out')
// (11, 10, 'neigh_op_bot_3')
// (12, 8, 'neigh_op_tnl_3')
// (12, 9, 'local_g1_3')
// (12, 9, 'lutff_6/in_0')
// (12, 9, 'neigh_op_lft_3')
// (12, 10, 'neigh_op_bnl_3')

reg n544 = 0;
// (10, 8, 'neigh_op_tnr_4')
// (10, 9, 'neigh_op_rgt_4')
// (10, 10, 'neigh_op_bnr_4')
// (11, 8, 'neigh_op_top_4')
// (11, 9, 'local_g1_4')
// (11, 9, 'lutff_4/out')
// (11, 9, 'lutff_5/in_0')
// (11, 10, 'neigh_op_bot_4')
// (12, 8, 'neigh_op_tnl_4')
// (12, 9, 'neigh_op_lft_4')
// (12, 10, 'neigh_op_bnl_4')

reg n545 = 0;
// (10, 8, 'neigh_op_tnr_6')
// (10, 9, 'neigh_op_rgt_6')
// (10, 10, 'neigh_op_bnr_6')
// (11, 8, 'neigh_op_top_6')
// (11, 9, 'local_g0_6')
// (11, 9, 'lutff_1/in_1')
// (11, 9, 'lutff_6/out')
// (11, 10, 'neigh_op_bot_6')
// (12, 8, 'neigh_op_tnl_6')
// (12, 9, 'neigh_op_lft_6')
// (12, 10, 'neigh_op_bnl_6')

wire \d_out[0] ;
// (10, 9, 'neigh_op_tnr_1')
// (10, 9, 'sp4_r_v_b_47')
// (10, 10, 'neigh_op_rgt_1')
// (10, 10, 'sp4_r_v_b_34')
// (10, 11, 'neigh_op_bnr_1')
// (10, 11, 'sp4_r_v_b_23')
// (10, 12, 'sp4_r_v_b_10')
// (11, 8, 'sp4_v_t_47')
// (11, 9, 'neigh_op_top_1')
// (11, 9, 'sp4_v_b_47')
// (11, 10, 'lutff_1/out')
// (11, 10, 'sp4_v_b_34')
// (11, 11, 'neigh_op_bot_1')
// (11, 11, 'sp4_v_b_23')
// (11, 12, 'sp4_h_r_4')
// (11, 12, 'sp4_v_b_10')
// (12, 9, 'neigh_op_tnl_1')
// (12, 10, 'neigh_op_lft_1')
// (12, 11, 'neigh_op_bnl_1')
// (12, 12, 'sp4_h_r_17')
// (13, 12, 'io_1/D_OUT_0')
// (13, 12, 'io_1/PAD')
// (13, 12, 'local_g0_1')
// (13, 12, 'span4_horz_17')

reg n547 = 0;
// (10, 9, 'neigh_op_tnr_2')
// (10, 10, 'neigh_op_rgt_2')
// (10, 11, 'neigh_op_bnr_2')
// (11, 9, 'neigh_op_top_2')
// (11, 10, 'local_g0_2')
// (11, 10, 'lutff_1/in_1')
// (11, 10, 'lutff_2/out')
// (11, 11, 'neigh_op_bot_2')
// (12, 9, 'neigh_op_tnl_2')
// (12, 10, 'neigh_op_lft_2')
// (12, 11, 'neigh_op_bnl_2')

reg n548 = 0;
// (10, 9, 'neigh_op_tnr_3')
// (10, 10, 'neigh_op_rgt_3')
// (10, 11, 'neigh_op_bnr_3')
// (11, 9, 'neigh_op_top_3')
// (11, 10, 'local_g1_3')
// (11, 10, 'lutff_3/out')
// (11, 10, 'lutff_6/in_0')
// (11, 11, 'neigh_op_bot_3')
// (12, 9, 'neigh_op_tnl_3')
// (12, 10, 'neigh_op_lft_3')
// (12, 11, 'neigh_op_bnl_3')

wire \d_out[1] ;
// (10, 10, 'neigh_op_tnr_1')
// (10, 11, 'neigh_op_rgt_1')
// (10, 12, 'neigh_op_bnr_1')
// (11, 9, 'sp4_r_v_b_43')
// (11, 10, 'neigh_op_top_1')
// (11, 10, 'sp4_r_v_b_30')
// (11, 11, 'lutff_1/out')
// (11, 11, 'sp4_r_v_b_19')
// (11, 12, 'neigh_op_bot_1')
// (11, 12, 'sp4_r_v_b_6')
// (12, 8, 'sp4_v_t_43')
// (12, 9, 'sp4_v_b_43')
// (12, 10, 'neigh_op_tnl_1')
// (12, 10, 'sp4_v_b_30')
// (12, 11, 'neigh_op_lft_1')
// (12, 11, 'sp4_v_b_19')
// (12, 12, 'neigh_op_bnl_1')
// (12, 12, 'sp4_h_r_0')
// (12, 12, 'sp4_v_b_6')
// (13, 12, 'io_0/D_OUT_0')
// (13, 12, 'io_0/PAD')
// (13, 12, 'local_g0_0')
// (13, 12, 'span4_horz_0')

reg n550 = 0;
// (10, 10, 'neigh_op_tnr_4')
// (10, 11, 'neigh_op_rgt_4')
// (10, 12, 'neigh_op_bnr_4')
// (11, 10, 'neigh_op_top_4')
// (11, 11, 'local_g0_4')
// (11, 11, 'lutff_1/in_1')
// (11, 11, 'lutff_4/out')
// (11, 12, 'neigh_op_bot_4')
// (12, 10, 'neigh_op_tnl_4')
// (12, 11, 'neigh_op_lft_4')
// (12, 12, 'neigh_op_bnl_4')

reg n551 = 0;
// (10, 10, 'neigh_op_tnr_7')
// (10, 11, 'neigh_op_rgt_7')
// (10, 12, 'neigh_op_bnr_7')
// (11, 10, 'neigh_op_top_7')
// (11, 11, 'local_g1_7')
// (11, 11, 'lutff_3/in_1')
// (11, 11, 'lutff_7/out')
// (11, 12, 'neigh_op_bot_7')
// (12, 10, 'neigh_op_tnl_7')
// (12, 11, 'neigh_op_lft_7')
// (12, 12, 'neigh_op_bnl_7')

reg n552 = 0;
// (10, 11, 'neigh_op_tnr_3')
// (10, 12, 'neigh_op_rgt_3')
// (10, 13, 'neigh_op_bnr_3')
// (11, 11, 'neigh_op_top_3')
// (11, 12, 'local_g1_3')
// (11, 12, 'lutff_2/in_0')
// (11, 12, 'lutff_3/out')
// (11, 13, 'neigh_op_bot_3')
// (12, 11, 'neigh_op_tnl_3')
// (12, 12, 'neigh_op_lft_3')
// (12, 13, 'neigh_op_bnl_3')

reg n553 = 0;
// (11, 5, 'neigh_op_tnr_4')
// (11, 6, 'neigh_op_rgt_4')
// (11, 7, 'neigh_op_bnr_4')
// (12, 5, 'neigh_op_top_4')
// (12, 6, 'local_g0_4')
// (12, 6, 'lutff_4/out')
// (12, 6, 'lutff_6/in_0')
// (12, 7, 'neigh_op_bot_4')
// (13, 5, 'logic_op_tnl_4')
// (13, 6, 'logic_op_lft_4')
// (13, 7, 'logic_op_bnl_4')

reg n554 = 0;
// (11, 5, 'neigh_op_tnr_5')
// (11, 6, 'neigh_op_rgt_5')
// (11, 7, 'neigh_op_bnr_5')
// (12, 5, 'neigh_op_top_5')
// (12, 6, 'local_g1_5')
// (12, 6, 'lutff_4/in_0')
// (12, 6, 'lutff_5/out')
// (12, 7, 'neigh_op_bot_5')
// (13, 5, 'logic_op_tnl_5')
// (13, 6, 'logic_op_lft_5')
// (13, 7, 'logic_op_bnl_5')

reg n555 = 0;
// (11, 6, 'neigh_op_tnr_0')
// (11, 7, 'neigh_op_rgt_0')
// (11, 8, 'neigh_op_bnr_0')
// (12, 6, 'local_g1_0')
// (12, 6, 'lutff_5/in_0')
// (12, 6, 'neigh_op_top_0')
// (12, 7, 'lutff_0/out')
// (12, 8, 'neigh_op_bot_0')
// (13, 6, 'logic_op_tnl_0')
// (13, 7, 'logic_op_lft_0')
// (13, 8, 'logic_op_bnl_0')

reg n556 = 0;
// (11, 6, 'neigh_op_tnr_2')
// (11, 7, 'neigh_op_rgt_2')
// (11, 8, 'neigh_op_bnr_2')
// (12, 6, 'neigh_op_top_2')
// (12, 7, 'local_g0_2')
// (12, 7, 'lutff_0/in_0')
// (12, 7, 'lutff_2/out')
// (12, 8, 'neigh_op_bot_2')
// (13, 6, 'logic_op_tnl_2')
// (13, 7, 'logic_op_lft_2')
// (13, 8, 'logic_op_bnl_2')

reg n557 = 0;
// (11, 8, 'neigh_op_tnr_5')
// (11, 9, 'neigh_op_rgt_5')
// (11, 10, 'neigh_op_bnr_5')
// (12, 8, 'neigh_op_top_5')
// (12, 9, 'local_g1_5')
// (12, 9, 'lutff_2/in_0')
// (12, 9, 'lutff_5/out')
// (12, 10, 'neigh_op_bot_5')
// (13, 8, 'logic_op_tnl_5')
// (13, 9, 'logic_op_lft_5')
// (13, 10, 'logic_op_bnl_5')

reg n558 = 0;
// (11, 8, 'neigh_op_tnr_6')
// (11, 9, 'neigh_op_rgt_6')
// (11, 10, 'neigh_op_bnr_6')
// (12, 8, 'neigh_op_top_6')
// (12, 9, 'local_g1_6')
// (12, 9, 'lutff_5/in_0')
// (12, 9, 'lutff_6/out')
// (12, 10, 'neigh_op_bot_6')
// (13, 8, 'logic_op_tnl_6')
// (13, 9, 'logic_op_lft_6')
// (13, 10, 'logic_op_bnl_6')

wire n559;
// (4, 3, 'lutff_0/cout')

wire n560;
// (2, 5, 'lutff_0/cout')

wire n561;
// (5, 12, 'lutff_6/lout')

wire n562;
// (9, 12, 'lutff_1/lout')

wire n563;
// (6, 8, 'lutff_4/lout')

wire n564;
// (5, 4, 'lutff_2/lout')

wire n565;
// (4, 8, 'lutff_5/lout')

wire n566;
// (7, 4, 'lutff_4/lout')

wire n567;
// (8, 8, 'lutff_6/lout')

wire n568;
// (7, 13, 'lutff_0/lout')

wire n569;
// (12, 6, 'lutff_5/lout')

wire n570;
// (5, 5, 'lutff_3/lout')

wire n571;
// (6, 12, 'lutff_1/lout')

wire n572;
// (7, 5, 'lutff_5/lout')

wire n573;
// (9, 5, 'lutff_7/lout')

wire n574;
// (6, 4, 'lutff_6/lout')

wire n575;
// (5, 9, 'lutff_0/lout')

wire n576;
// (7, 9, 'lutff_2/lout')

wire n577;
// (9, 9, 'lutff_4/lout')

wire n578;
// (5, 8, 'lutff_4/lout')

wire n579;
// (7, 8, 'lutff_6/lout')

wire n580;
// (2, 7, 'lutff_6/lout')

wire n581;
// (6, 11, 'lutff_5/lout')

wire n582;
// (8, 11, 'lutff_7/lout')

wire n583;
// (5, 12, 'lutff_1/lout')

wire n584;
// (7, 12, 'lutff_3/lout')

wire n585;
// (4, 8, 'lutff_0/lout')

wire n586;
// (9, 12, 'lutff_5/lout')

wire n587;
// (2, 8, 'lutff_7/lout')

wire n588;
// (8, 8, 'lutff_1/lout')

wire n589;
// (2, 11, 'lutff_3/lout')

wire n590;
// (11, 10, 'lutff_2/lout')

wire n591;
// (7, 13, 'lutff_4/lout')

wire n592;
// (7, 5, 'lutff_0/lout')

wire n593;
// (12, 9, 'lutff_5/lout')

wire n594;
// (5, 5, 'lutff_7/lout')

wire n595;
// (9, 5, 'lutff_2/lout')

wire n596;
// (4, 12, 'lutff_6/lout')

wire n597;
// (8, 4, 'lutff_3/lout')

wire n598;
// (6, 15, 'lutff_7/lout')

wire n599;
// (6, 7, 'lutff_3/lout')

wire n600;
// (8, 7, 'lutff_5/lout')

wire n601;
// (7, 8, 'lutff_1/lout')

wire n602;
// (9, 8, 'lutff_3/lout')

wire n603;
// (5, 11, 'lutff_4/lout')

wire n604;
// (7, 11, 'lutff_6/lout')

wire n605;
// (6, 11, 'lutff_0/lout')

wire n606;
// (11, 9, 'lutff_5/lout')

wire n607;
// (5, 12, 'lutff_5/lout')

wire n608;
// (9, 12, 'lutff_0/lout')

wire n609;
// (2, 8, 'lutff_2/lout')

wire n610;
// (5, 4, 'lutff_1/lout')

wire n611;
// (6, 8, 'lutff_3/lout')

wire n612;
// (4, 8, 'lutff_4/lout')

wire n613;
// (7, 4, 'lutff_3/lout')

wire n614;
// (8, 8, 'lutff_5/lout')

wire n615;
// (7, 12, 'lutff_7/lout')

wire n616;
// (11, 10, 'lutff_6/lout')

wire n617;
// (6, 3, 'lutff_1/lout')

wire n618;
// (6, 14, 'lutff_1/lout')

wire n619;
// (8, 3, 'lutff_3/lout')

wire n620;
// (6, 6, 'lutff_6/lout')

wire n621;
// (4, 11, 'lutff_5/lout')

wire n622;
// (8, 7, 'lutff_0/lout')

wire n623;
// (6, 7, 'lutff_7/lout')

wire n624;
// (11, 5, 'lutff_3/lout')

wire n625;
// (5, 8, 'lutff_3/lout')

wire n626;
// (7, 11, 'lutff_1/lout')

wire n627;
// (4, 7, 'lutff_7/lout')

wire n628;
// (6, 11, 'lutff_4/lout')

wire n629;
// (8, 11, 'lutff_6/lout')

wire n630;
// (5, 12, 'lutff_0/lout')

wire n631;
// (5, 4, 'lutff_5/lout')

wire n632;
// (2, 11, 'lutff_2/lout')

wire n633;
// (7, 4, 'lutff_7/lout')

wire n634;
// (11, 10, 'lutff_1/lout')

wire n635;
// (6, 3, 'lutff_5/lout')

wire n636;
// (6, 14, 'lutff_5/lout')

wire n637;
// (8, 3, 'lutff_7/lout')

wire n638;
// (7, 15, 'lutff_3/lout')

wire n639;
// (9, 4, 'lutff_5/lout')

wire n640;
// (5, 7, 'lutff_6/lout')

wire n641;
// (6, 7, 'lutff_2/lout')

wire n642;
// (8, 7, 'lutff_4/lout')

wire n643;
// (11, 5, 'lutff_7/lout')

wire n644;
// (7, 8, 'lutff_0/lout')

wire n645;
// (5, 8, 'lutff_7/lout')

wire n646;
// (2, 7, 'lutff_0/lout')

wire n647;
// (7, 11, 'lutff_5/lout')

wire n648;
// (4, 7, 'lutff_2/lout')

wire n649;
// (8, 11, 'lutff_1/lout')

wire n650;
// (6, 10, 'lutff_3/lout')

wire n651;
// (11, 9, 'lutff_4/lout')

wire n652;
// (8, 10, 'lutff_5/lout')

wire n653;
// (7, 4, 'lutff_2/lout')

wire n654;
// (7, 3, 'lutff_6/lout')

wire n655;
// (4, 10, 'lutff_3/lout')

wire n656;
// (6, 14, 'lutff_0/lout')

wire n657;
// (6, 3, 'lutff_0/lout')

wire n658;
// (8, 3, 'lutff_2/lout')

wire n659;
// (2, 2, 'lutff_6/lout')

wire n660;
// (9, 4, 'lutff_0/lout')

wire n661;
// (5, 7, 'lutff_1/lout')

wire n662;
// (7, 15, 'lutff_7/lout')

wire n663;
// (4, 11, 'lutff_4/lout')

wire n664;
// (7, 7, 'lutff_3/lout')

wire n665;
// (6, 15, 'lutff_1/lout')

wire n666;
// (4, 3, 'lutff_0/out')

wire n667;
// (4, 3, 'lutff_0/lout')

wire n668;
// (4, 3, 'carry_in_mux')

// Carry-In for (4 3)
assign n668 = 1;

wire n669;
// (9, 7, 'lutff_5/lout')

wire n670;
// (5, 8, 'lutff_2/lout')

wire n671;
// (7, 8, 'lutff_4/lout')

wire n672;
// (7, 11, 'lutff_0/lout')

wire n673;
// (9, 8, 'lutff_6/lout')

wire n674;
// (5, 11, 'lutff_7/lout')

wire n675;
// (2, 7, 'lutff_4/lout')

wire n676;
// (4, 7, 'lutff_6/lout')

wire n677;
// (11, 6, 'lutff_3/lout')

wire n678;
// (8, 10, 'lutff_0/lout')

wire n679;
// (6, 10, 'lutff_7/lout')

wire n680;
// (6, 13, 'lutff_3/lout')

wire n681;
// (6, 2, 'lutff_3/lout')

wire n682;
// (8, 2, 'lutff_5/lout')

wire n683;
// (7, 3, 'lutff_1/lout')

wire n684;
// (5, 6, 'lutff_4/lout')

wire n685;
// (4, 10, 'lutff_7/lout')

wire n686;
// (6, 3, 'lutff_4/lout')

wire n687;
// (6, 14, 'lutff_4/lout')

wire n688;
// (4, 2, 'lutff_3/lout')

wire n689;
// (8, 3, 'lutff_6/lout')

wire n690;
// (7, 15, 'lutff_2/lout')

wire n691;
// (5, 7, 'lutff_5/lout')

wire n692;
// (9, 7, 'lutff_0/lout')

wire n693;
// (7, 7, 'lutff_7/lout')

wire n694;
// (4, 3, 'lutff_4/lout')

wire n695;
// (11, 5, 'lutff_6/lout')

wire n696;
// (6, 9, 'lutff_1/lout')

wire n697;
// (8, 6, 'lutff_7/lout')

wire n698;
// (2, 6, 'lutff_3/lout')

wire n699;
// (5, 14, 'lutff_4/lout')

wire n700;
// (12, 7, 'lutff_2/lout')

wire n701;
// (6, 10, 'lutff_2/lout')

wire n702;
// (8, 10, 'lutff_4/lout')

wire n703;
// (8, 2, 'lutff_0/lout')

wire n704;
// (6, 13, 'lutff_7/lout')

wire n705;
// (6, 2, 'lutff_7/lout')

wire n706;
// (9, 11, 'lutff_2/lout')

wire n707;
// (5, 3, 'lutff_3/lout')

wire n708;
// (7, 3, 'lutff_5/lout')

wire n709;
// (4, 10, 'lutff_2/lout')

wire n710;
// (9, 3, 'lutff_7/lout')

wire n711;
// (8, 3, 'lutff_1/lout')

wire n712;
// (4, 2, 'lutff_7/lout')

wire n713;
// (5, 7, 'lutff_0/lout')

wire n714;
// (9, 7, 'lutff_4/lout')

wire n715;
// (5, 10, 'lutff_2/lout')

wire n716;
// (7, 10, 'lutff_4/lout')

wire n717;
// (11, 5, 'lutff_1/lout')

wire n718;
// (8, 6, 'lutff_2/lout')

wire n719;
// (5, 13, 'lutff_7/lout')

wire n720;
// (2, 9, 'lutff_4/lout')

wire n721;
// (6, 9, 'lutff_5/lout')

wire n722;
// (8, 9, 'lutff_7/lout')

wire n723;
// (4, 6, 'lutff_0/lout')

wire n724;
// (2, 6, 'lutff_7/lout')

wire n725;
// (5, 2, 'lutff_6/lout')

wire n726;
// (6, 10, 'lutff_6/lout')

wire n727;
// (6, 13, 'lutff_2/lout')

wire n728;
// (6, 2, 'lutff_2/lout')

wire n729;
// (7, 3, 'lutff_0/lout')

wire n730;
// (5, 6, 'lutff_3/lout')

wire n731;
// (4, 10, 'lutff_6/lout')

wire n732;
// (4, 2, 'lutff_2/lout')

wire n733;
// (8, 13, 'lutff_0/lout')

wire n734;
// (6, 5, 'lutff_3/lout')

wire n735;
// (8, 5, 'lutff_5/lout')

wire n736;
// (5, 10, 'lutff_6/lout')

wire n737;
// (9, 10, 'lutff_1/lout')

wire n738;
// (5, 13, 'lutff_2/lout')

wire n739;
// (7, 2, 'lutff_4/lout')

wire n740;
// (8, 6, 'lutff_6/lout')

wire n741;
// (4, 9, 'lutff_1/lout')

wire n742;
// (8, 9, 'lutff_2/lout')

wire n743;
// (5, 14, 'lutff_3/lout')

wire n744;
// (6, 10, 'lutff_1/lout')

wire n745;
// (7, 14, 'lutff_5/lout')

wire n746;
// (8, 10, 'lutff_3/lout')

wire n747;
// (6, 2, 'lutff_6/lout')

wire n748;
// (6, 13, 'lutff_6/lout')

wire n749;
// (9, 11, 'lutff_1/lout')

wire n750;
// (7, 3, 'lutff_4/lout')

wire n751;
// (4, 10, 'lutff_1/lout')

wire n752;
// (5, 6, 'lutff_7/lout')

wire n753;
// (2, 2, 'lutff_4/lout')

wire n754;
// (4, 2, 'lutff_6/lout')

wire n755;
// (7, 6, 'lutff_6/lout')

wire n756;
// (4, 13, 'lutff_3/lout')

wire n757;
// (8, 13, 'lutff_4/lout')

wire n758;
// (11, 12, 'lutff_3/lout')

wire n759;
// (8, 5, 'lutff_0/lout')

wire n760;
// (2, 5, 'lutff_6/lout')

wire n761;
// (6, 5, 'lutff_7/lout')

wire n762;
// (11, 11, 'lutff_7/lout')

wire n763;
// (5, 10, 'lutff_1/lout')

wire n764;
// (7, 10, 'lutff_3/lout')

wire n765;
// (8, 6, 'lutff_1/lout')

wire n766;
// (9, 10, 'lutff_5/lout')

wire n767;
// (5, 13, 'lutff_6/lout')

wire n768;
// (2, 9, 'lutff_3/lout')

wire n769;
// (6, 9, 'lutff_4/lout')

wire n770;
// (4, 9, 'lutff_5/lout')

wire n771;
// (8, 9, 'lutff_6/lout')

wire n772;
// (11, 7, 'lutff_0/lout')

wire n773;
// (7, 14, 'lutff_0/lout')

wire n774;
// (5, 2, 'lutff_5/lout')

wire n775;
// (11, 8, 'lutff_1/lout')

wire n776;
// (6, 12, 'lutff_5/lout')

wire n777;
// (6, 4, 'lutff_1/lout')

wire n778;
// (2, 13, 'lutff_5/lout')

wire n779;
// (5, 9, 'lutff_4/lout')

wire n780;
// (4, 13, 'lutff_7/lout')

wire n781;
// (6, 5, 'lutff_2/lout')

wire n782;
// (7, 9, 'lutff_6/lout')

wire n783;
// (2, 5, 'lutff_1/out')

wire n784;
// (2, 5, 'lutff_1/lout')

wire n785;
// (8, 5, 'lutff_4/lout')

wire n786;
// (9, 10, 'lutff_0/lout')

wire n787;
// (7, 10, 'lutff_7/lout')

wire n788;
// (5, 13, 'lutff_1/lout')

wire n789;
// (7, 2, 'lutff_3/lout')

wire n790;
// (8, 9, 'lutff_1/lout')

wire n791;
// (2, 9, 'lutff_7/lout')

wire n792;
// (11, 7, 'lutff_4/lout')

wire n793;
// (12, 7, 'lutff_0/lout')

wire n794;
// (4, 6, 'lutff_3/lout')

wire n795;
// (12, 6, 'lutff_4/lout')

wire n796;
// (5, 5, 'lutff_2/lout')

wire n797;
// (7, 5, 'lutff_4/lout')

wire n798;
// (6, 12, 'lutff_0/lout')

wire n799;
// (4, 12, 'lutff_1/lout')

wire n800;
// (9, 5, 'lutff_6/lout')

wire n801;
// (8, 12, 'lutff_2/lout')

wire n802;
// (2, 4, 'lutff_4/lout')

wire n803;
// (6, 4, 'lutff_5/lout')

wire n804;
// (8, 4, 'lutff_7/lout')

wire n805;
// (2, 13, 'lutff_0/lout')

wire n806;
// (7, 9, 'lutff_1/lout')

wire n807;
// (9, 6, 'lutff_7/lout')

wire n808;
// (9, 9, 'lutff_3/lout')

wire n809;
// (2, 5, 'lutff_5/lout')

wire n810;
// (6, 5, 'lutff_6/lout')

wire n811;
// (7, 10, 'lutff_2/lout')

wire n812;
// (9, 10, 'lutff_4/lout')

wire n813;
// (5, 13, 'lutff_5/lout')

wire n814;
// (2, 9, 'lutff_2/lout')

wire n815;
// (7, 2, 'lutff_7/lout')

wire n816;
// (4, 9, 'lutff_4/lout')

wire n817;
// (8, 8, 'lutff_0/lout')

wire n818;
// (6, 8, 'lutff_7/lout')

wire n819;
// (9, 13, 'lutff_5/lout')

wire n820;
// (9, 5, 'lutff_1/lout')

wire n821;
// (6, 4, 'lutff_0/lout')

wire n822;
// (8, 12, 'lutff_6/lout')

wire n823;
// (8, 4, 'lutff_2/lout')

wire n824;
// (9, 6, 'lutff_2/lout')

wire n825;
// (2, 13, 'lutff_4/lout')

wire n826;
// (2, 5, 'lutff_0/out')

wire n827;
// (2, 5, 'lutff_0/lout')

wire n828;
// (2, 5, 'carry_in_mux')

// Carry-In for (2 5)
assign n828 = 1;

wire n829;
// (4, 13, 'lutff_6/lout')

wire n830;
// (6, 5, 'lutff_1/lout')

wire n831;
// (7, 9, 'lutff_5/lout')

wire n832;
// (11, 11, 'lutff_1/lout')

wire n833;
// (8, 5, 'lutff_3/lout')

wire n834;
// (9, 9, 'lutff_7/lout')

wire n835;
// (5, 12, 'lutff_4/lout')

wire n836;
// (7, 12, 'lutff_6/lout')

wire n837;
// (11, 7, 'lutff_3/lout')

wire n838;
// (4, 8, 'lutff_3/lout')

wire n839;
// (2, 11, 'lutff_6/lout')

wire n840;
// (7, 13, 'lutff_7/lout')

wire n841;
// (7, 5, 'lutff_3/lout')

wire n842;
// (9, 5, 'lutff_5/lout')

wire n843;
// (2, 12, 'lutff_7/lout')

wire n844;
// (8, 12, 'lutff_1/lout')

wire n845;
// (2, 4, 'lutff_3/lout')

wire n846;
// (6, 4, 'lutff_4/lout')

wire n847;
// (8, 4, 'lutff_6/lout')

wire n848;
// (6, 7, 'lutff_6/lout')

wire n849;
// (7, 9, 'lutff_0/lout')

wire n850;
// (9, 9, 'lutff_2/lout')

wire n851;
// (6, 11, 'lutff_3/lout')

wire n852;
// (7, 12, 'lutff_1/lout')

wire n853;
// (9, 12, 'lutff_3/lout')

wire n854;
// (6, 8, 'lutff_6/lout')

wire n855;
// (2, 11, 'lutff_1/lout')

wire n856;
// (7, 4, 'lutff_6/lout')

wire n857;
// (4, 8, 'lutff_7/lout')

wire n858;
// (7, 5, 'lutff_7/lout')

wire n859;
// (4, 12, 'lutff_4/lout')

wire n860;
// (8, 4, 'lutff_1/lout')

wire n861;
// (6, 15, 'lutff_5/lout')

wire n862;
// (6, 7, 'lutff_1/lout')

wire n863;
// (8, 7, 'lutff_3/lout')

wire n864;
// (5, 8, 'lutff_6/lout')

wire n865;
// (9, 8, 'lutff_1/lout')

wire n866;
// (5, 11, 'lutff_2/lout')

wire n867;
// (7, 11, 'lutff_4/lout')

wire n868;
// (4, 7, 'lutff_1/lout')

wire n869;
// (8, 11, 'lutff_0/lout')

wire n870;
// (6, 11, 'lutff_7/lout')

wire n871;
// (11, 9, 'lutff_3/lout')

wire n872;
// (5, 12, 'lutff_3/lout')

wire n873;
// (7, 12, 'lutff_5/lout')

wire n874;
// (4, 8, 'lutff_2/lout')

wire n875;
// (7, 4, 'lutff_1/lout')

wire n876;
// (2, 11, 'lutff_5/lout')

wire n877;
// (11, 10, 'lutff_4/lout')

wire n878;
// (7, 5, 'lutff_2/lout')

wire n879;
// (9, 5, 'lutff_4/lout')

wire n880;
// (2, 4, 'lutff_2/lout')

wire n881;
// (4, 11, 'lutff_3/lout')

wire n882;
// (6, 15, 'lutff_0/lout')

wire n883;
// (6, 7, 'lutff_5/lout')

wire n884;
// (11, 13, 'lutff_5/lout')

wire n885;
// (8, 7, 'lutff_7/lout')

wire n886;
// (5, 8, 'lutff_1/lout')

wire n887;
// (7, 8, 'lutff_3/lout')

wire n888;
// (9, 8, 'lutff_5/lout')

wire n889;
// (5, 11, 'lutff_6/lout')

wire n890;
// (4, 7, 'lutff_5/lout')

wire n891;
// (6, 11, 'lutff_2/lout')

wire n892;
// (11, 6, 'lutff_2/lout')

wire n893;
// (8, 11, 'lutff_4/lout')

wire n894;
// (11, 9, 'lutff_7/lout')

wire n895;
// (7, 12, 'lutff_0/lout')

wire n896;
// (5, 12, 'lutff_7/lout')

wire n897;
// (4, 8, 'lutff_6/lout')

wire n898;
// (7, 4, 'lutff_5/lout')

wire n899;
// (2, 11, 'lutff_0/lout')

wire n900;
// (6, 14, 'lutff_3/lout')

wire n901;
// (6, 3, 'lutff_3/lout')

wire n902;
// (8, 3, 'lutff_5/lout')

wire n903;
// (12, 9, 'lutff_2/lout')

wire n904;
// (7, 15, 'lutff_1/lout')

wire n905;
// (9, 4, 'lutff_3/lout')

wire n906;
// (5, 7, 'lutff_4/lout')

wire n907;
// (6, 15, 'lutff_4/lout')

wire n908;
// (4, 3, 'lutff_3/lout')

wire n909;
// (6, 7, 'lutff_0/lout')

wire n910;
// (8, 7, 'lutff_2/lout')

wire n911;
// (11, 5, 'lutff_5/lout')

wire n912;
// (5, 8, 'lutff_5/lout')

wire n913;
// (9, 8, 'lutff_0/lout')

wire n914;
// (7, 8, 'lutff_7/lout')

wire n915;
// (5, 11, 'lutff_1/lout')

wire n916;
// (7, 11, 'lutff_3/lout')

wire n917;
// (4, 7, 'lutff_0/lout')

wire n918;
// (2, 7, 'lutff_7/lout')

wire n919;
// (11, 6, 'lutff_6/lout')

wire n920;
// (5, 12, 'lutff_2/lout')

wire n921;
// (7, 12, 'lutff_4/lout')

wire n922;
// (4, 8, 'lutff_1/lout')

wire n923;
// (7, 4, 'lutff_0/lout')

wire n924;
// (9, 12, 'lutff_6/lout')

wire n925;
// (8, 3, 'lutff_0/lout')

wire n926;
// (6, 3, 'lutff_7/lout')

wire n927;
// (6, 6, 'lutff_3/lout')

wire n928;
// (7, 15, 'lutff_5/lout')

wire n929;
// (4, 11, 'lutff_2/lout')

wire n930;
// (9, 4, 'lutff_7/lout')

wire n931;
// (9, 7, 'lutff_3/lout')

wire n932;
// (2, 14, 'lutff_5/lout')

wire n933;
// (6, 7, 'lutff_4/lout')

wire n934;
// (8, 7, 'lutff_6/lout')

wire n935;
// (11, 5, 'lutff_0/lout')

wire n936;
// (5, 8, 'lutff_0/lout')

wire n937;
// (7, 8, 'lutff_2/lout')

wire n938;
// (7, 11, 'lutff_7/lout')

wire n939;
// (5, 14, 'lutff_7/lout')

wire n940;
// (6, 10, 'lutff_5/lout')

wire n941;
// (11, 9, 'lutff_6/lout')

wire n942;
// (6, 2, 'lutff_1/lout')

wire n943;
// (6, 13, 'lutff_1/lout')

wire n944;
// (8, 2, 'lutff_3/lout')

wire n945;
// (9, 11, 'lutff_5/lout')

wire n946;
// (5, 6, 'lutff_2/lout')

wire n947;
// (4, 10, 'lutff_5/lout')

wire n948;
// (6, 3, 'lutff_2/lout')

wire n949;
// (6, 14, 'lutff_2/lout')

wire n950;
// (4, 2, 'lutff_1/lout')

wire n951;
// (8, 3, 'lutff_4/lout')

wire n952;
// (7, 15, 'lutff_0/lout')

wire n953;
// (5, 7, 'lutff_3/lout')

wire n954;
// (7, 7, 'lutff_5/lout')

wire n955;
// (4, 3, 'lutff_2/lout')

wire n956;
// (9, 7, 'lutff_7/lout')

wire n957;
// (8, 7, 'lutff_1/lout')

wire n958;
// (8, 6, 'lutff_5/lout')

wire n959;
// (7, 11, 'lutff_2/lout')

wire n960;
// (2, 6, 'lutff_1/lout')

wire n961;
// (6, 10, 'lutff_0/lout')

wire n962;
// (11, 9, 'lutff_1/lout')

wire n963;
// (8, 10, 'lutff_2/lout')

wire n964;
// (6, 2, 'lutff_5/lout')

wire n965;
// (8, 2, 'lutff_7/lout')

wire n966;
// (7, 3, 'lutff_3/lout')

wire n967;
// (4, 10, 'lutff_0/lout')

wire n968;
// (2, 10, 'lutff_7/lout')

wire n969;
// (5, 6, 'lutff_6/lout')

wire n970;
// (6, 3, 'lutff_6/lout')

wire n971;
// (6, 14, 'lutff_6/lout')

wire n972;
// (4, 2, 'lutff_5/lout')

wire n973;
// (11, 12, 'lutff_2/lout')

wire n974;
// (11, 4, 'lutff_7/lout')

wire n975;
// (4, 11, 'lutff_1/lout')

wire n976;
// (7, 7, 'lutff_0/lout')

wire n977;
// (9, 4, 'lutff_6/lout')

wire n978;
// (5, 7, 'lutff_7/lout')

wire n979;
// (9, 7, 'lutff_2/lout')

wire n980;
// (4, 3, 'lutff_6/lout')

wire n981;
// (4, 14, 'lutff_6/lout')

wire n982;
// (8, 6, 'lutff_0/lout')

wire n983;
// (6, 9, 'lutff_3/lout')

wire n984;
// (5, 2, 'lutff_4/lout')

wire n985;
// (4, 6, 'lutff_7/lout')

wire n986;
// (6, 10, 'lutff_4/lout')

wire n987;
// (6, 13, 'lutff_0/lout')

wire n988;
// (8, 10, 'lutff_6/lout')

wire n989;
// (2, 10, 'lutff_2/lout')

wire n990;
// (5, 6, 'lutff_1/lout')

wire n991;
// (7, 3, 'lutff_7/lout')

wire n992;
// (4, 10, 'lutff_4/lout')

wire n993;
// (4, 2, 'lutff_0/lout')

wire n994;
// (8, 13, 'lutff_7/lout')

wire n995;
// (11, 4, 'lutff_2/lout')

wire n996;
// (5, 7, 'lutff_2/lout')

wire n997;
// (4, 3, 'lutff_1/out')

wire n998;
// (4, 3, 'lutff_1/lout')

wire n999;
// (9, 7, 'lutff_6/lout')

wire n1000;
// (5, 13, 'lutff_0/lout')

wire n1001;
// (7, 10, 'lutff_6/lout')

wire n1002;
// (7, 2, 'lutff_2/lout')

wire n1003;
// (8, 6, 'lutff_4/lout')

wire n1004;
// (8, 9, 'lutff_0/lout')

wire n1005;
// (6, 9, 'lutff_7/lout')

wire n1006;
// (2, 6, 'lutff_0/lout')

wire n1007;
// (5, 14, 'lutff_1/lout')

wire n1008;
// (4, 6, 'lutff_2/lout')

wire n1009;
// (7, 14, 'lutff_3/lout')

wire n1010;
// (8, 10, 'lutff_1/lout')

wire n1011;
// (6, 13, 'lutff_4/lout')

wire n1012;
// (8, 2, 'lutff_6/lout')

wire n1013;
// (7, 3, 'lutff_2/lout')

wire n1014;
// (5, 6, 'lutff_5/lout')

wire n1015;
// (4, 2, 'lutff_4/lout')

wire n1016;
// (5, 9, 'lutff_7/lout')

wire n1017;
// (2, 5, 'lutff_4/lout')

wire n1018;
// (6, 5, 'lutff_5/lout')

wire n1019;
// (11, 4, 'lutff_6/lout')

wire n1020;
// (8, 5, 'lutff_7/lout')

wire n1021;
// (7, 10, 'lutff_1/lout')

wire n1022;
// (9, 10, 'lutff_3/lout')

wire n1023;
// (6, 9, 'lutff_2/lout')

wire n1024;
// (7, 2, 'lutff_6/lout')

wire n1025;
// (4, 9, 'lutff_3/lout')

wire n1026;
// (8, 9, 'lutff_4/lout')

wire n1027;
// (5, 2, 'lutff_3/lout')

wire n1028;
// (5, 14, 'lutff_5/lout')

wire n1029;
// (4, 6, 'lutff_6/lout')

wire n1030;
// (7, 14, 'lutff_7/lout')

wire n1031;
// (8, 2, 'lutff_1/lout')

wire n1032;
// (6, 12, 'lutff_3/lout')

wire n1033;
// (8, 12, 'lutff_5/lout')

wire n1034;
// (5, 6, 'lutff_0/lout')

wire n1035;
// (9, 6, 'lutff_1/lout')

wire n1036;
// (2, 13, 'lutff_3/lout')

wire n1037;
// (5, 9, 'lutff_2/lout')

wire n1038;
// (4, 13, 'lutff_5/lout')

wire n1039;
// (7, 9, 'lutff_4/lout')

wire n1040;
// (8, 5, 'lutff_2/lout')

wire n1041;
// (9, 9, 'lutff_6/lout')

wire n1042;
// (11, 3, 'lutff_5/lout')

wire n1043;
// (7, 10, 'lutff_5/lout')

wire n1044;
// (7, 2, 'lutff_1/lout')

wire n1045;
// (8, 6, 'lutff_3/lout')

wire n1046;
// (9, 10, 'lutff_7/lout')

wire n1047;
// (6, 9, 'lutff_6/lout')

wire n1048;
// (4, 6, 'lutff_1/lout')

wire n1049;
// (5, 2, 'lutff_7/lout')

wire n1050;
// (11, 8, 'lutff_3/lout')

wire n1051;
// (8, 12, 'lutff_0/lout')

wire n1052;
// (6, 12, 'lutff_7/lout')

wire n1053;
// (6, 4, 'lutff_3/lout')

wire n1054;
// (8, 4, 'lutff_5/lout')

wire n1055;
// (4, 13, 'lutff_0/lout')

wire n1056;
// (8, 13, 'lutff_1/lout')

wire n1057;
// (2, 13, 'lutff_7/lout')

wire n1058;
// (9, 6, 'lutff_5/lout')

wire n1059;
// (5, 9, 'lutff_6/lout')

wire n1060;
// (2, 5, 'lutff_3/lout')

wire n1061;
// (6, 5, 'lutff_4/lout')

wire n1062;
// (9, 9, 'lutff_1/lout')

wire n1063;
// (4, 5, 'lutff_5/lout')

wire n1064;
// (8, 5, 'lutff_6/lout')

wire n1065;
// (11, 11, 'lutff_4/lout')

wire n1066;
// (7, 10, 'lutff_0/lout')

wire n1067;
// (5, 10, 'lutff_7/lout')

wire n1068;
// (9, 10, 'lutff_2/lout')

wire n1069;
// (5, 13, 'lutff_3/lout')

wire n1070;
// (4, 9, 'lutff_2/lout')

wire n1071;
// (8, 9, 'lutff_3/lout')

wire n1072;
// (6, 8, 'lutff_5/lout')

wire n1073;
// (8, 8, 'lutff_7/lout')

wire n1074;
// (5, 2, 'lutff_2/lout')

wire n1075;
// (7, 13, 'lutff_1/lout')

wire n1076;
// (12, 6, 'lutff_6/lout')

wire n1077;
// (5, 5, 'lutff_4/lout')

wire n1078;
// (7, 5, 'lutff_6/lout')

wire n1079;
// (6, 12, 'lutff_2/lout')

wire n1080;
// (4, 12, 'lutff_3/lout')

wire n1081;
// (8, 12, 'lutff_4/lout')

wire n1082;
// (1, 8, 'lutff_6/lout')

wire n1083;
// (8, 4, 'lutff_0/lout')

wire n1084;
// (6, 4, 'lutff_7/lout')

wire n1085;
// (9, 6, 'lutff_0/lout')

wire n1086;
// (2, 13, 'lutff_2/lout')

wire n1087;
// (7, 6, 'lutff_7/lout')

wire n1088;
// (4, 13, 'lutff_4/lout')

wire n1089;
// (7, 9, 'lutff_3/lout')

wire n1090;
// (8, 13, 'lutff_5/lout')

wire n1091;
// (8, 5, 'lutff_1/lout')

wire n1092;
// (2, 5, 'lutff_7/lout')

wire n1093;
// (9, 9, 'lutff_5/lout')

wire n1094;
// (6, 11, 'lutff_6/lout')

wire n1095;
// (7, 2, 'lutff_0/lout')

wire n1096;
// (6, 8, 'lutff_0/lout')

wire n1097;
// (11, 7, 'lutff_1/lout')

wire n1098;
// (8, 8, 'lutff_2/lout')

wire n1099;
// (11, 10, 'lutff_3/lout')

wire n1100;
// (7, 13, 'lutff_5/lout')

wire n1101;
// (12, 9, 'lutff_6/lout')

wire n1102;
// (9, 5, 'lutff_3/lout')

wire n1103;
// (6, 12, 'lutff_6/lout')

wire n1104;
// (2, 4, 'lutff_1/lout')

wire n1105;
// (6, 4, 'lutff_2/lout')

wire n1106;
// (4, 12, 'lutff_7/lout')

wire n1107;
// (8, 4, 'lutff_4/lout')

wire n1108;
// (7, 6, 'lutff_2/lout')

wire n1109;
// (9, 6, 'lutff_4/lout')

wire n1110;
// (5, 9, 'lutff_5/lout')

wire n1111;
// (9, 9, 'lutff_0/lout')

wire n1112;
// (2, 5, 'lutff_2/lout')

wire n1113;
// (7, 9, 'lutff_7/lout')

wire n1114;
// (4, 5, 'lutff_4/lout')

wire n1115;
// (11, 11, 'lutff_3/lout')

wire n1116;
// (6, 11, 'lutff_1/lout')

wire n1117;
// (8, 11, 'lutff_3/lout')

assign n667  = /* LUT    4  3  0 */ 1'b0;
assign n784  = /* LUT    2  5  1 */ 1'b0;
assign n827  = /* LUT    2  5  0 */ 1'b0;
assign n998  = /* LUT    4  3  1 */ 1'b0;
assign n561  = /* LUT    5 12  6 */ (n202 ? n34 : (n102 ? n147 : !n147));
assign n562  = /* LUT    9 12  1 */ n530;
assign n563  = /* LUT    6  8  4 */ n24;
assign n564  = /* LUT    5  4  2 */ (n51 ? 1'b0 : !n52);
assign n565  = /* LUT    4  8  5 */ (n190 ? (n188 ? (n132 ? !n133 : n133) : (n132 ? n133 : !n133)) : (n188 ? (n132 ? n133 : !n133) : (n132 ? !n133 : n133)));
assign n566  = /* LUT    7  4  4 */ (n168 ? (n329 ? (n250 ? !n336 : n336) : (n250 ? n336 : !n336)) : 1'b0);
assign n567  = /* LUT    8  8  6 */ n448;
assign n568  = /* LUT    7 13  0 */ (n387 ? (n59 ? (n60 ? !n397 : 1'b1) : 1'b1) : 1'b0);
assign n569  = /* LUT   12  6  5 */ n555;
assign n570  = /* LUT    5  5  3 */ n261;
assign n571  = /* LUT    6 12  1 */ (n59 ? (n60 ? 1'b1 : !n109) : (n60 ? !n301 : 1'b1));
assign n572  = /* LUT    7  5  5 */ (n431 ? (n257 ? (n332 ? 1'b1 : !n168) : (n332 ? !n168 : 1'b1)) : (n257 ? (n332 ? 1'b0 : n168) : (n332 ? n168 : 1'b0)));
assign n573  = /* LUT    9  5  7 */ n392;
assign n574  = /* LUT    6  4  6 */ (n13 ? n91 : 1'b0);
assign n575  = /* LUT    5  9  0 */ (n281 ? (n216 ? (n263 ? n212 : !n212) : (n263 ? !n212 : n212)) : (n216 ? (n263 ? !n212 : n212) : (n263 ? n212 : !n212)));
assign n576  = /* LUT    7  9  2 */ (n376 ? (n59 ? (n60 ? !n30 : 1'b1) : 1'b1) : 1'b0);
assign n577  = /* LUT    9  9  4 */ n455;
assign n578  = /* LUT    5  8  4 */ (n195 ? (n185 ? (n198 ? n133 : !n133) : (n198 ? !n133 : n133)) : (n185 ? (n198 ? !n133 : n133) : (n198 ? n133 : !n133)));
assign n579  = /* LUT    7  8  6 */ (n21 ? n357 : n360);
assign n580  = /* LUT    2  7  6 */ n57;
assign n581  = /* LUT    6 11  5 */ (n21 ? n295 : n293);
assign n582  = /* LUT    8 11  7 */ (n59 ? (n60 ? n474 : n461) : n474);
assign n583  = /* LUT    5 12  1 */ (n162 ? (n59 ? (n60 ? !n34 : 1'b1) : 1'b1) : 1'b0);
assign n584  = /* LUT    7 12  3 */ n298;
assign n585  = /* LUT    4  8  0 */ (n194 ? n132 : !n132);
assign n586  = /* LUT    9 12  5 */ n392;
assign n587  = /* LUT    2  8  7 */ !n57;
assign n588  = /* LUT    8  8  1 */ n449;
assign n589  = /* LUT    2 11  3 */ n77;
assign n590  = /* LUT   11 10  2 */ (n196 ? n423 : !n423);
assign n591  = /* LUT    7 13  4 */ (n59 ? (n60 ? 1'b1 : !n303) : (n60 ? !n110 : 1'b1));
assign n592  = /* LUT    7  5  0 */ (n4 ? !n259 : 1'b0);
assign n593  = /* LUT   12  9  5 */ n558;
assign n594  = /* LUT    5  5  7 */ (n104 ? !n255 : n255);
assign n595  = /* LUT    9  5  2 */ (n490 ? !n507 : !n494);
assign n596  = /* LUT    4 12  6 */ n159;
assign n597  = /* LUT    8  4  3 */ (n406 ? !n418 : n418);
assign n598  = /* LUT    6 15  7 */ (n59 ? (n60 ? n310 : n318) : n310);
assign n599  = /* LUT    6  7  3 */ (n200 ? (n178 ? n144 : !n144) : 1'b0);
assign n600  = /* LUT    8  7  5 */ n497;
assign n601  = /* LUT    7  8  1 */ (n22 ? n25 : !n25);
assign n602  = /* LUT    9  8  3 */ n423;
assign n603  = /* LUT    5 11  4 */ n220;
assign n604  = /* LUT    7 11  6 */ n214;
assign n605  = /* LUT    6 11  0 */ (n21 ? !n292 : !n294);
assign n606  = /* LUT   11  9  5 */ n544;
assign n607  = /* LUT    5 12  5 */ n158;
assign n608  = /* LUT    9 12  0 */ n533;
assign n609  = /* LUT    2  8  2 */ (n22 ? (n62 ? !n65 : 1'b1) : (n62 ? n65 : 1'b0));
assign n610  = /* LUT    5  4  1 */ (n11 ? (n41 ? 1'b1 : (n6 ? 1'b1 : n92)) : 1'b0);
assign n611  = /* LUT    6  8  3 */ (n269 ? (n197 ? (n62 ? n356 : 1'b0) : (n62 ? !n356 : 1'b1)) : (n197 ? (n62 ? !n356 : 1'b1) : (n62 ? n356 : 1'b0)));
assign n612  = /* LUT    4  8  4 */ (n188 ? (n194 ? (n132 ? n133 : !n133) : (n132 ? !n133 : n133)) : (n194 ? (n132 ? !n133 : n133) : (n132 ? n133 : !n133)));
assign n613  = /* LUT    7  4  3 */ (n177 ? (n340 ? (n173 ? !n337 : n337) : (n173 ? n337 : !n337)) : (n340 ? (n173 ? n337 : !n337) : (n173 ? !n337 : n337)));
assign n614  = /* LUT    8  8  5 */ (n458 ? (n446 ? n169 : 1'b1) : (n446 ? !n169 : 1'b0));
assign n615  = /* LUT    7 12  7 */ n384;
assign n616  = /* LUT   11 10  6 */ n548;
assign n617  = /* LUT    6  3  1 */ (n325 ? (n324 ? n239 : (n239 ? 1'b0 : !n87)) : (n324 ? n239 : (n239 ? 1'b1 : n87)));
assign n618  = /* LUT    6 14  1 */ (n311 ? (n59 ? (n60 ? !n318 : 1'b1) : 1'b1) : 1'b0);
assign n619  = /* LUT    8  3  3 */ (n424 ? !n418 : n418);
assign n620  = /* LUT    6  6  6 */ (n197 ? !n346 : n346);
assign n621  = /* LUT    4 11  5 */ (n104 ? (n62 ? !n155 : 1'b1) : (n62 ? n155 : 1'b0));
assign n622  = /* LUT    8  7  0 */ (n470 ? (n423 ? n169 : 1'b1) : (n423 ? !n169 : 1'b0));
assign n623  = /* LUT    6  7  7 */ n255;
assign n624  = /* LUT   11  5  3 */ (n537 ? (n41 ? 1'b1 : (n6 ? 1'b1 : n92)) : 1'b0);
assign n625  = /* LUT    5  8  3 */ (n189 ? (n266 ? (n270 ? !n205 : n205) : !n270) : (n266 ? n205 : 1'b0));
assign n626  = /* LUT    7 11  1 */ n381;
assign n627  = /* LUT    4  7  7 */ (n54 ? (n130 ? (n128 ? !n131 : n131) : (n128 ? n131 : 1'b0)) : (n130 ? (n128 ? 1'b0 : !n131) : 1'b1));
assign n628  = /* LUT    6 11  4 */ (n140 ? (n62 ? !n292 : 1'b1) : (n62 ? n292 : 1'b0));
assign n629  = /* LUT    8 11  6 */ n469;
assign n630  = /* LUT    5 12  0 */ (n226 ? (n90 ? (n153 ? !n202 : 1'b1) : (n153 ? 1'b1 : !n202)) : 1'b0);
assign n631  = /* LUT    5  4  5 */ (n51 ? (n14 ? (n50 ? 1'b0 : !n52) : 1'b0) : 1'b0);
assign n632  = /* LUT    2 11  2 */ n75;
assign n633  = /* LUT    7  4  7 */ (n351 ? (n41 ? 1'b1 : (n6 ? 1'b1 : n92)) : 1'b0);
assign n634  = /* LUT   11 10  1 */ (select ? n423 : n547);
assign n635  = /* LUT    6  3  5 */ (n324 ? n238 : (n239 ? n325 : 1'b1));
assign n636  = /* LUT    6 14  5 */ (n59 ? (n60 ? n303 : n312) : n303);
assign n637  = /* LUT    8  3  7 */ (n416 ? (n406 ? !n418 : n418) : (n406 ? n418 : !n418));
assign n638  = /* LUT    7 15  3 */ (n59 ? (n60 ? n400 : n397) : n400);
assign n639  = /* LUT    9  4  5 */ (n500 ? (n41 ? 1'b0 : (n6 ? 1'b0 : !n92)) : 1'b0);
assign n640  = /* LUT    5  7  6 */ (n180 ? (n200 ? n263 : 1'b1) : (n200 ? (n263 ? n187 : !n187) : !n187));
assign n641  = /* LUT    6  7  2 */ (n103 ? (n7 ? n201 : !n201) : (n7 ? !n201 : n201));
assign n642  = /* LUT    8  7  4 */ n439;
assign n643  = /* LUT   11  5  7 */ n534;
assign n644  = /* LUT    7  8  0 */ (n21 ? !n356 : !n359);
assign n645  = /* LUT    5  8  7 */ n23;
assign n646  = /* LUT    2  7  0 */ (n55 ? n17 : 1'b0);
assign n647  = /* LUT    7 11  5 */ n347;
assign n648  = /* LUT    4  7  2 */ (n186 ? (n63 ? (n135 ? n136 : !n136) : n135) : (n63 ? 1'b1 : n136));
assign n649  = /* LUT    8 11  1 */ n471;
assign n650  = /* LUT    6 10  3 */ (n21 ? n288 : n207);
assign n651  = /* LUT   11  9  4 */ n70;
assign n652  = /* LUT    8 10  5 */ n464;
assign n653  = /* LUT    7  4  2 */ (n333 ? (n340 ? (n173 ? n334 : !n334) : (n173 ? !n334 : n334)) : (n340 ? (n173 ? !n334 : n334) : (n173 ? n334 : !n334)));
assign n654  = /* LUT    7  3  6 */ (n236 ? (n254 ? !n88 : 1'b1) : (n254 ? n88 : 1'b0));
assign n655  = /* LUT    4 10  3 */ (n197 ? (n62 ? !n28 : 1'b1) : (n62 ? n28 : 1'b0));
assign n656  = /* LUT    6 14  0 */ (n59 ? (n60 ? 1'b1 : !n310) : (n60 ? !n111 : 1'b1));
assign n657  = /* LUT    6  3  0 */ (n324 ? (n325 ? n87 : (n87 ? 1'b0 : !n239)) : (n325 ? n87 : (n87 ? 1'b1 : n239)));
assign n658  = /* LUT    8  3  2 */ (n419 ? (n404 ? (n485 ? n413 : !n413) : n485) : (n404 ? 1'b0 : n413));
assign n659  = /* LUT    2  2  6 */ (n8 ? (n42 ? !rst : 1'b0) : 1'b0);
assign n660  = /* LUT    9  4  0 */ (n409 ? (n176 ? 1'b1 : n495) : (n176 ? n487 : (n495 ? n487 : !n487)));
assign n661  = /* LUT    5  7  1 */ (n263 ? (n200 ? !n180 : 1'b0) : (n200 ? (n180 ? n268 : !n268) : !n268));
assign n662  = /* LUT    7 15  7 */ n399;
assign n663  = /* LUT    4 11  4 */ (n21 ? n155 : n154);
assign n664  = /* LUT    7  7  3 */ n353;
assign n665  = /* LUT    6 15  1 */ n316;
assign n669  = /* LUT    9  7  5 */ n504;
assign n670  = /* LUT    5  8  2 */ (n205 ? (n266 ? (n189 ? n191 : !n191) : n191) : (n266 ? n189 : 1'b0));
assign n671  = /* LUT    7  8  4 */ (n22 ? (n271 ? (n23 ? n62 : 1'b0) : (n23 ? !n62 : 1'b1)) : (n271 ? (n23 ? !n62 : 1'b1) : (n23 ? n62 : 1'b0)));
assign n672  = /* LUT    7 11  0 */ (n59 ? (n60 ? 1'b1 : !n224) : (n60 ? !n379 : 1'b1));
assign n673  = /* LUT    9  8  6 */ n446;
assign n674  = /* LUT    5 11  7 */ n76;
assign n675  = /* LUT    2  7  4 */ (n55 ? (n17 ? 1'b1 : n49) : (n17 ? n49 : 1'b1));
assign n676  = /* LUT    4  7  6 */ (n128 ? (n54 ? (n130 ? !n131 : 1'b0) : (n130 ? n131 : !n131)) : (n54 ? (n130 ? n131 : 1'b1) : n131));
assign n677  = /* LUT   11  6  3 */ n460;
assign n678  = /* LUT    8 10  0 */ n466;
assign n679  = /* LUT    6 10  7 */ (n25 ? (n62 ? n286 : 1'b0) : (n62 ? !n286 : 1'b1));
assign n680  = /* LUT    6 13  3 */ (n202 ? n318 : (n137 ? n282 : !n282));
assign n681  = /* LUT    6  2  3 */ (n87 ? (n327 ? (n240 ? !n326 : n326) : (n240 ? n326 : !n326)) : 1'b0);
assign n682  = /* LUT    8  2  5 */ (n484 ? n407 : !n407);
assign n683  = /* LUT    7  3  1 */ (n237 ? (n173 ? (n88 ? n248 : 1'b1) : (n88 ? !n248 : 1'b0)) : (n173 ? (n88 ? !n248 : 1'b0) : (n88 ? n248 : 1'b1)));
assign n684  = /* LUT    5  6  4 */ (n178 ? (n184 ? (n263 ? n186 : !n186) : n263) : (n184 ? n186 : 1'b1));
assign n685  = /* LUT    4 10  7 */ (n21 ? n28 : n68);
assign n686  = /* LUT    6  3  4 */ (n237 ? (n242 ? 1'b1 : n243) : (n242 ? 1'b0 : !n243));
assign n687  = /* LUT    6 14  4 */ n313;
assign n688  = /* LUT    4  2  3 */ (n122 ? (n123 ? (n120 ? 1'b0 : !n121) : 1'b0) : 1'b0);
assign n689  = /* LUT    8  3  6 */ (n9 ? (n413 ? !n342 : n342) : 1'b0);
assign n690  = /* LUT    7 15  2 */ n394;
assign n691  = /* LUT    5  7  5 */ (n203 ? n107 : !n107);
assign n692  = /* LUT    9  7  0 */ (n498 ? (n142 ? n169 : 1'b1) : (n142 ? !n169 : 1'b0));
assign n693  = /* LUT    7  7  7 */ n352;
assign n694  = /* LUT    4  3  4 */ (n122 ? 1'b0 : (n168 ? (n58 ? 1'b1 : n8) : 1'b1));
assign n695  = /* LUT   11  5  6 */ n535;
assign n696  = /* LUT    6  9  1 */ (n21 ? !n280 : !n276);
assign n697  = /* LUT    8  6  7 */ n432;
assign n698  = /* LUT    2  6  3 */ (n101 ? (n16 ? n18 : !n18) : (n16 ? !n18 : n18));
assign n699  = /* LUT    5 14  4 */ (n59 ? (n60 ? n228 : n225) : n228);
assign n700  = /* LUT   12  7  2 */ n539;
assign n701  = /* LUT    6 10  2 */ n213;
assign n702  = /* LUT    8 10  4 */ n468;
assign n703  = /* LUT    8  2  0 */ (n484 ? (n407 ? n404 : !n404) : (n407 ? !n404 : n404));
assign n704  = /* LUT    6 13  7 */ n33;
assign n705  = /* LUT    6  2  7 */ (n242 ? n248 : !n248);
assign n706  = /* LUT    9 11  2 */ n525;
assign n707  = /* LUT    5  3  3 */ (n8 ? 1'b0 : (n41 ? 1'b0 : (n6 ? 1'b0 : !n4)));
assign n708  = /* LUT    7  3  5 */ (n411 ? (n331 ? (n328 ? !n245 : n245) : (n328 ? n245 : !n245)) : (n331 ? (n328 ? n245 : !n245) : (n328 ? !n245 : n245)));
assign n709  = /* LUT    4 10  2 */ (n138 ? (n146 ? (n29 ? !n62 : 1'b1) : (n29 ? n62 : 1'b0)) : (n146 ? (n29 ? n62 : 1'b0) : (n29 ? !n62 : 1'b1)));
assign n710  = /* LUT    9  3  7 */ (n485 ? (n406 ? !n418 : n418) : (n406 ? n418 : !n418));
assign n711  = /* LUT    8  3  1 */ (n404 ? (n485 ? (n419 ? !n413 : n413) : !n413) : (n485 ? 1'b1 : !n419));
assign n712  = /* LUT    4  2  7 */ (rst ? 1'b0 : (n6 ? 1'b1 : (n41 ? !n113 : 1'b0)));
assign n713  = /* LUT    5  7  0 */ (n103 ? (n201 ? n205 : !n205) : (n201 ? !n205 : n205));
assign n714  = /* LUT    9  7  4 */ n511;
assign n715  = /* LUT    5 10  2 */ n215;
assign n716  = /* LUT    7 10  4 */ (n21 ? n370 : n373);
assign n717  = /* LUT   11  5  1 */ (n538 ? (n41 ? 1'b1 : (n6 ? 1'b1 : n92)) : 1'b0);
assign n718  = /* LUT    8  6  2 */ n434;
assign n719  = /* LUT    5 13  7 */ (n60 ? (n59 ? n230 : n225) : n230);
assign n720  = /* LUT    2  9  4 */ (n21 ? n71 : n67);
assign n721  = /* LUT    6  9  5 */ (n104 ? (n62 ? !n280 : 1'b1) : (n62 ? n280 : 1'b0));
assign n722  = /* LUT    8  9  7 */ n467;
assign n723  = /* LUT    4  6  0 */ (n182 ? (n129 ? (n186 ? n184 : 1'b1) : (n186 ? !n184 : 1'b0)) : (n129 ? (n186 ? !n184 : 1'b0) : (n186 ? n184 : 1'b1)));
assign n724  = /* LUT    2  6  7 */ (n17 ? !n55 : n55);
assign n725  = /* LUT    5  2  6 */ (rst ? 1'b0 : (n166 ? 1'b1 : (n41 ? n113 : 1'b0)));
assign n726  = /* LUT    6 10  6 */ (n368 ? (n289 ? !n62 : 1'b1) : (n289 ? n62 : 1'b0));
assign n727  = /* LUT    6 13  2 */ (n59 ? (n60 ? n109 : n307) : n109);
assign n728  = /* LUT    6  2  2 */ (n241 ? 1'b0 : (n322 ? 1'b0 : (n325 ? n238 : 1'b1)));
assign n729  = /* LUT    7  3  0 */ (n402 ? (n408 ? 1'b1 : n246) : (n408 ? n247 : (n246 ? n247 : !n247)));
assign n730  = /* LUT    5  6  3 */ (n178 ? !n201 : n201);
assign n731  = /* LUT    4 10  6 */ (n21 ? n148 : n152);
assign n732  = /* LUT    4  2  2 */ (n2 ? (n58 ? 1'b1 : rst) : 1'b1);
assign n733  = /* LUT    8 13  0 */ n482;
assign n734  = /* LUT    6  5  3 */ (n4 ? (n252 ? (n14 ? !n52 : n52) : 1'b0) : 1'b0);
assign n735  = /* LUT    8  5  5 */ (n437 ? 1'b0 : !n425);
assign n736  = /* LUT    5 10  6 */ n289;
assign n737  = /* LUT    9 10  1 */ n519;
assign n738  = /* LUT    5 13  2 */ n36;
assign n739  = /* LUT    7  2  4 */ (n323 ? n321 : !n321);
assign n740  = /* LUT    8  6  6 */ n427;
assign n741  = /* LUT    4  9  1 */ (n104 ? n138 : !n138);
assign n742  = /* LUT    8  9  2 */ n457;
assign n743  = /* LUT    5 14  3 */ n233;
assign n744  = /* LUT    6 10  1 */ (n196 ? (n62 ? n288 : 1'b0) : (n62 ? !n288 : 1'b1));
assign n745  = /* LUT    7 14  5 */ n393;
assign n746  = /* LUT    8 10  3 */ n380;
assign n747  = /* LUT    6  2  6 */ (n242 ? (n248 ? 1'b0 : !n320) : (n248 ? !n320 : 1'b0));
assign n748  = /* LUT    6 13  6 */ n305;
assign n749  = /* LUT    9 11  1 */ n531;
assign n750  = /* LUT    7  3  4 */ (n89 ? (n407 ? n246 : 1'b1) : (n407 ? (n246 ? n247 : !n247) : n247));
assign n751  = /* LUT    4 10  1 */ (n21 ? !n145 : !n151);
assign n752  = /* LUT    5  6  7 */ (n107 ? (n178 ? (n201 ? !n205 : n205) : (n201 ? n205 : !n205)) : (n178 ? (n201 ? n205 : !n205) : (n201 ? !n205 : n205)));
assign n753  = /* LUT    2  2  4 */ (rst ? 1'b0 : (n4 ? 1'b1 : (n8 ? !n42 : 1'b0)));
assign n754  = /* LUT    4  2  6 */ (n122 ? (n123 ? (n120 ? n121 : 1'b0) : 1'b0) : 1'b0);
assign n755  = /* LUT    7  6  6 */ n428;
assign n756  = /* LUT    4 13  3 */ n165;
assign n757  = /* LUT    8 13  4 */ n483;
assign n758  = /* LUT   11 12  3 */ n529;
assign n759  = /* LUT    8  5  0 */ (n429 ? (n343 ? (n344 ? 1'b1 : !n168) : (n344 ? !n168 : 1'b1)) : (n343 ? (n344 ? 1'b0 : n168) : (n344 ? n168 : 1'b0)));
assign n760  = /* LUT    2  5  6 */ (n97 ? !n52 : n52);
assign n761  = /* LUT    6  5  7 */ n179;
assign n762  = /* LUT   11 11  7 */ (n271 ? !n421 : n421);
assign n763  = /* LUT    5 10  1 */ n149;
assign n764  = /* LUT    7 10  3 */ (n140 ? (n62 ? !n372 : 1'b1) : (n62 ? n372 : 1'b0));
assign n765  = /* LUT    8  6  1 */ n435;
assign n766  = /* LUT    9 10  5 */ n517;
assign n767  = /* LUT    5 13  6 */ n218;
assign n768  = /* LUT    2  9  3 */ (n105 ? (n62 ? !n71 : 1'b1) : (n62 ? n71 : 1'b0));
assign n769  = /* LUT    6  9  4 */ (n25 ? (n62 ? n275 : 1'b0) : (n62 ? !n275 : 1'b1));
assign n770  = /* LUT    4  9  5 */ (n139 ? !n25 : n25);
assign n771  = /* LUT    8  9  6 */ (n463 ? (n262 ? n169 : 1'b1) : (n262 ? !n169 : 1'b0));
assign n772  = /* LUT   11  7  0 */ n541;
assign n773  = /* LUT    7 14  0 */ (n59 ? (n60 ? 1'b1 : !n400) : (n60 ? !n395 : 1'b1));
assign n774  = /* LUT    5  2  5 */ (rst ? 1'b1 : (n58 ? !n118 : 1'b0));
assign n775  = /* LUT   11  8  1 */ n459;
assign n776  = /* LUT    6 12  5 */ n302;
assign n777  = /* LUT    6  4  1 */ (n337 ? (n245 ? (n249 ? n252 : 1'b1) : (n249 ? !n252 : 1'b0)) : (n245 ? (n249 ? !n252 : 1'b0) : (n249 ? n252 : 1'b1)));
assign n778  = /* LUT    2 13  5 */ n80;
assign n779  = /* LUT    5  9  4 */ (n103 ? n216 : !n216);
assign n780  = /* LUT    4 13  7 */ n163;
assign n781  = /* LUT    6  5  2 */ (n4 ? (n260 ? (n51 ? !n50 : 1'b0) : 1'b0) : 1'b0);
assign n782  = /* LUT    7  9  6 */ (n202 ? n30 : (n460 ? n354 : !n354));
assign n785  = /* LUT    8  5  4 */ (n434 ? (n41 ? 1'b0 : (n6 ? 1'b0 : !n92)) : 1'b0);
assign n786  = /* LUT    9 10  0 */ n524;
assign n787  = /* LUT    7 10  7 */ (n21 ? n372 : n27);
assign n788  = /* LUT    5 13  1 */ (n59 ? (n60 ? 1'b1 : !n228) : (n60 ? !n230 : 1'b1));
assign n789  = /* LUT    7  2  3 */ (n403 ? (n242 ? (n248 ? 1'b0 : !n320) : (n248 ? !n320 : 1'b0)) : (n242 ? (n248 ? 1'b1 : n320) : (n248 ? n320 : 1'b1)));
assign n790  = /* LUT    8  9  1 */ (n59 ? (n60 ? 1'b1 : !n474) : (n60 ? !n26 : 1'b1));
assign n791  = /* LUT    2  9  7 */ (n21 ? n72 : n69);
assign n792  = /* LUT   11  7  4 */ n540;
assign n793  = /* LUT   12  7  0 */ n556;
assign n794  = /* LUT    4  6  3 */ (n18 ? (n129 ? !n183 : n183) : (n129 ? n183 : !n183));
assign n795  = /* LUT   12  6  4 */ n554;
assign n796  = /* LUT    5  5  2 */ (select ? n255 : n175);
assign n797  = /* LUT    7  5  4 */ (n353 ? (n41 ? 1'b0 : (n6 ? 1'b0 : !n92)) : 1'b0);
assign n798  = /* LUT    6 12  0 */ (n84 ? (n59 ? (n60 ? !n307 : 1'b1) : 1'b1) : 1'b0);
assign n799  = /* LUT    4 12  1 */ n31;
assign n800  = /* LUT    9  5  6 */ (n426 ? 1'b0 : !n492);
assign n801  = /* LUT    8 12  2 */ n475;
assign n802  = /* LUT    2  4  4 */ n90;
assign n803  = /* LUT    6  4  5 */ (n4 ? (n14 ? 1'b1 : n50) : 1'b0);
assign n804  = /* LUT    8  4  7 */ (n489 ? (n10 ? (n417 ? !n168 : 1'b1) : (n417 ? 1'b1 : !n168)) : (n10 ? (n417 ? n168 : 1'b0) : (n417 ? 1'b0 : n168)));
assign n805  = /* LUT    2 13  0 */ (n60 ? (n59 ? n37 : n34) : n37);
assign n806  = /* LUT    7  9  1 */ (n452 ? (n428 ? (n274 ? !n202 : 1'b1) : (n274 ? 1'b1 : !n202)) : 1'b0);
assign n807  = /* LUT    9  6  7 */ n512;
assign n808  = /* LUT    9  9  3 */ n374;
assign n809  = /* LUT    2  5  5 */ (n96 ? !n51 : n51);
assign n810  = /* LUT    6  5  6 */ (n52 ? !n14 : 1'b0);
assign n811  = /* LUT    7 10  2 */ (n140 ? (n62 ? !n370 : 1'b1) : (n62 ? n370 : 1'b0));
assign n812  = /* LUT    9 10  4 */ n518;
assign n813  = /* LUT    5 13  5 */ n231;
assign n814  = /* LUT    2  9  2 */ (n21 ? !n65 : !n66);
assign n815  = /* LUT    7  2  7 */ (n242 ? (n402 ? n89 : 1'b0) : (n410 ? (n402 ? n89 : 1'b0) : (n402 ? !n89 : 1'b1)));
assign n816  = /* LUT    4  9  4 */ (n105 ? (n62 ? !n72 : 1'b1) : (n62 ? n72 : 1'b0));
assign n817  = /* LUT    8  8  0 */ (n450 ? !n339 : n339);
assign n818  = /* LUT    6  8  7 */ n272;
assign n819  = /* LUT    9 13  5 */ n421;
assign n820  = /* LUT    9  5  1 */ (n41 ? 1'b0 : (n6 ? 1'b0 : !n92));
assign n821  = /* LUT    6  4  0 */ (n13 ? (n52 ? 1'b0 : (n51 ? !n14 : 1'b1)) : 1'b0);
assign n822  = /* LUT    8 12  6 */ n478;
assign n823  = /* LUT    8  4  2 */ (n126 ? (n409 ? 1'b0 : !n487) : (n409 ? !n345 : (n487 ? !n345 : n345)));
assign n824  = /* LUT    9  6  2 */ n500;
assign n825  = /* LUT    2 13  4 */ n81;
assign n829  = /* LUT    4 13  6 */ n164;
assign n830  = /* LUT    6  5  1 */ (n265 ? (n256 ? (n338 ? 1'b1 : !n168) : (n338 ? !n168 : 1'b1)) : (n256 ? (n338 ? 1'b0 : n168) : (n338 ? n168 : 1'b0)));
assign n831  = /* LUT    7  9  5 */ n363;
assign n832  = /* LUT   11 11  1 */ (select ? n262 : n550);
assign n833  = /* LUT    8  5  3 */ (n437 ? (n499 ? 1'b1 : n422) : (n499 ? n425 : (n422 ? n425 : !n425)));
assign n834  = /* LUT    9  9  7 */ n515;
assign n835  = /* LUT    5 12  4 */ n221;
assign n836  = /* LUT    7 12  6 */ n386;
assign n837  = /* LUT   11  7  3 */ n102;
assign n838  = /* LUT    4  8  3 */ (n134 ? (n195 ? (n138 ? n141 : !n141) : (n138 ? !n141 : n141)) : (n195 ? (n138 ? !n141 : n141) : (n138 ? n141 : !n141)));
assign n839  = /* LUT    2 11  6 */ n108;
assign n840  = /* LUT    7 13  7 */ (n202 ? n312 : (n347 ? n367 : !n367));
assign n841  = /* LUT    7  5  3 */ (n336 ? (n330 ? !n332 : n332) : (n330 ? n332 : !n332));
assign n842  = /* LUT    9  5  5 */ (n524 ? (n41 ? 1'b0 : (n6 ? 1'b0 : !n92)) : 1'b0);
assign n843  = /* LUT    2 12  7 */ n85;
assign n844  = /* LUT    8 12  1 */ n479;
assign n845  = /* LUT    2  4  3 */ (n43 ? (n52 ? (n14 ? 1'b0 : !n50) : n14) : 1'b0);
assign n846  = /* LUT    6  4  4 */ (n50 ? !n51 : 1'b0);
assign n847  = /* LUT    8  4  6 */ (n126 ? 1'b0 : !n345);
assign n848  = /* LUT    6  7  6 */ (n131 ? (n128 ? (n130 ? n54 : 1'b1) : (n130 ? 1'b1 : n54)) : (n128 ? n54 : 1'b0));
assign n849  = /* LUT    7  9  0 */ (n202 ? (n460 ? n354 : !n354) : 1'b0);
assign n850  = /* LUT    9  9  2 */ n520;
assign n851  = /* LUT    6 11  3 */ (n21 ? n296 : n208);
assign n852  = /* LUT    7 12  1 */ n383;
assign n853  = /* LUT    9 12  3 */ n528;
assign n854  = /* LUT    6  8  6 */ (n284 ? (n255 ? n169 : 1'b1) : (n255 ? !n169 : 1'b0));
assign n855  = /* LUT    2 11  1 */ n73;
assign n856  = /* LUT    7  4  6 */ (n168 ? (n45 ? (n329 ? n336 : !n336) : (n329 ? !n336 : n336)) : 1'b0);
assign n857  = /* LUT    4  8  7 */ (n198 ? n133 : !n133);
assign n858  = /* LUT    7  5  7 */ n99;
assign n859  = /* LUT    4 12  4 */ n160;
assign n860  = /* LUT    8  4  1 */ (n488 ? (n485 ? !n420 : n420) : (n485 ? n420 : !n420));
assign n861  = /* LUT    6 15  5 */ n315;
assign n862  = /* LUT    6  7  1 */ (n54 ? (n131 ? 1'b0 : n128) : (n131 ? 1'b1 : n130));
assign n863  = /* LUT    8  7  3 */ n443;
assign n864  = /* LUT    5  8  6 */ (n193 ? (n266 ? !n201 : 1'b0) : (n266 ? (n201 ? !n191 : n191) : n191));
assign n865  = /* LUT    9  8  1 */ (select ? n446 : n451);
assign n866  = /* LUT    5 11  2 */ (n210 ? (n102 ? (n147 ? !n202 : 1'b1) : (n147 ? 1'b1 : !n202)) : 1'b0);
assign n867  = /* LUT    7 11  4 */ n364;
assign n868  = /* LUT    4  7  1 */ (n186 ? (n63 ? !n136 : (n135 ? !n136 : n136)) : (n63 ? 1'b0 : !n135));
assign n869  = /* LUT    8 11  0 */ n472;
assign n870  = /* LUT    6 11  7 */ (n271 ? (n140 ? (n290 ? n62 : 1'b0) : (n290 ? !n62 : 1'b1)) : (n140 ? (n290 ? !n62 : 1'b1) : (n290 ? n62 : 1'b0)));
assign n871  = /* LUT   11  9  3 */ n456;
assign n872  = /* LUT    5 12  3 */ n217;
assign n873  = /* LUT    7 12  5 */ (n202 ? n397 : (n392 ? n64 : !n64));
assign n874  = /* LUT    4  8  2 */ (n195 ? (n185 ? (n61 ? !n62 : 1'b1) : (n61 ? n62 : 1'b0)) : (n185 ? (n61 ? n62 : 1'b0) : (n61 ? !n62 : 1'b1)));
assign n875  = /* LUT    7  4  1 */ (n333 ? (n334 ? !n329 : n329) : (n334 ? n329 : !n329));
assign n876  = /* LUT    2 11  5 */ n74;
assign n877  = /* LUT   11 10  4 */ n522;
assign n878  = /* LUT    7  5  2 */ (n348 ? (n258 ? (n336 ? !n168 : 1'b1) : (n336 ? 1'b1 : !n168)) : (n258 ? (n336 ? n168 : 1'b0) : (n336 ? 1'b0 : n168)));
assign n879  = /* LUT    9  5  4 */ (n496 ? (n41 ? 1'b0 : (n6 ? 1'b0 : !n92)) : 1'b0);
assign n880  = /* LUT    2  4  2 */ (n50 ? (n14 ? n91 : 1'b0) : 1'b0);
assign n881  = /* LUT    4 11  3 */ (n104 ? (n62 ? !n150 : 1'b1) : (n62 ? n150 : 1'b0));
assign n882  = /* LUT    6 15  0 */ n319;
assign n883  = /* LUT    6  7  5 */ (n267 ? (n20 ? (n178 ? n268 : 1'b1) : (n178 ? !n268 : 1'b0)) : (n20 ? (n178 ? !n268 : 1'b0) : (n178 ? n268 : 1'b1)));
assign n884  = /* LUT   11 13  5 */ n32;
assign n885  = /* LUT    8  7  7 */ n506;
assign n886  = /* LUT    5  8  1 */ (n7 ? !n205 : n205);
assign n887  = /* LUT    7  8  3 */ (n355 ? (n62 ? !n358 : 1'b1) : (n62 ? n358 : 1'b0));
assign n888  = /* LUT    9  8  5 */ n142;
assign n889  = /* LUT    5 11  6 */ (n59 ? (n60 ? n224 : n30) : n224);
assign n890  = /* LUT    4  7  5 */ (n184 ? (n127 ? !n135 : 1'b0) : (n127 ? (n135 ? !n136 : n136) : !n136));
assign n891  = /* LUT    6 11  2 */ (n271 ? (n62 ? !n295 : 1'b1) : (n62 ? n295 : 1'b0));
assign n892  = /* LUT   11  6  2 */ n137;
assign n893  = /* LUT    8 11  4 */ n473;
assign n894  = /* LUT   11  9  7 */ n209;
assign n895  = /* LUT    7 12  0 */ (n388 ? (n392 ? (n64 ? !n202 : 1'b1) : (n64 ? 1'b1 : !n202)) : 1'b0);
assign n896  = /* LUT    5 12  7 */ (n202 ? n225 : (n90 ? n153 : !n153));
assign n897  = /* LUT    4  8  6 */ (n190 ? (n132 ? (n195 ? !n185 : n185) : (n195 ? n185 : !n185)) : (n132 ? (n195 ? n185 : !n185) : (n195 ? !n185 : n185)));
assign n898  = /* LUT    7  4  5 */ (n404 ? (n9 ? n419 : 1'b1) : (n9 ? (n419 ? n46 : !n46) : !n46));
assign n899  = /* LUT    2 11  0 */ n78;
assign n900  = /* LUT    6 14  3 */ (n60 ? (n59 ? n111 : n318) : n111);
assign n901  = /* LUT    6  3  3 */ (n87 ? (n239 ? n324 : (n325 ? n324 : 1'b1)) : (n239 ? 1'b0 : (n325 ? 1'b1 : n324)));
assign n902  = /* LUT    8  3  5 */ (n416 ? (n424 ? !n406 : n406) : (n424 ? n406 : !n406));
assign n903  = /* LUT   12  9  2 */ n557;
assign n904  = /* LUT    7 15  1 */ n396;
assign n905  = /* LUT    9  4  3 */ (n486 ? (n12 ? 1'b1 : n491) : (n12 ? 1'b0 : !n491));
assign n906  = /* LUT    5  7  4 */ (n144 ? (n200 ? n178 : 1'b0) : (n200 ? (n178 ? n187 : !n187) : n187));
assign n907  = /* LUT    6 15  4 */ n317;
assign n908  = /* LUT    4  3  3 */ (n171 ? (n121 ? 1'b0 : !n117) : (n121 ? !n117 : 1'b0));
assign n909  = /* LUT    6  7  0 */ (n130 ? (n128 ? !n131 : 1'b0) : (n128 ? n54 : 1'b1));
assign n910  = /* LUT    8  7  2 */ n441;
assign n911  = /* LUT   11  5  5 */ n444;
assign n912  = /* LUT    5  8  5 */ (n192 ? (n20 ? (n134 ? !n185 : n185) : (n134 ? n185 : !n185)) : (n20 ? (n134 ? n185 : !n185) : (n134 ? !n185 : n185)));
assign n913  = /* LUT    9  8  0 */ (n169 ? !n92 : 1'b0);
assign n914  = /* LUT    7  8  7 */ (n21 ? n358 : n199);
assign n915  = /* LUT    5 11  1 */ (n211 ? (n216 ? (n263 ? !n212 : n212) : (n263 ? n212 : !n212)) : (n216 ? (n263 ? n212 : !n212) : (n263 ? !n212 : n212)));
assign n916  = /* LUT    7 11  3 */ n377;
assign n917  = /* LUT    4  7  0 */ (n184 ? (n127 ? n136 : 1'b1) : (n135 ? (n127 ? 1'b1 : n136) : (n127 ? 1'b0 : !n136)));
assign n918  = /* LUT    2  7  7 */ (n17 ? 1'b1 : (n48 ? (n55 ? 1'b1 : n49) : 1'b0));
assign n919  = /* LUT   11  6  6 */ n102;
assign n920  = /* LUT    5 12  2 */ n222;
assign n921  = /* LUT    7 12  4 */ n382;
assign n922  = /* LUT    4  8  1 */ !n21;
assign n923  = /* LUT    7  4  0 */ (n419 ? (n9 ? !n404 : 1'b0) : (n9 ? (n404 ? n244 : !n244) : !n244));
assign n924  = /* LUT    9 12  6 */ n527;
assign n925  = /* LUT    8  3  0 */ (n413 ? (n9 ? n342 : 1'b1) : (n9 ? (n342 ? !n244 : n244) : n244));
assign n926  = /* LUT    6  3  7 */ (n325 ? (n324 ? (n87 ? n239 : !n239) : (n87 ? 1'b0 : n239)) : (n324 ? (n87 ? !n239 : 1'b0) : 1'b1));
assign n927  = /* LUT    6  6  3 */ (select ? n346 : n264);
assign n928  = /* LUT    7 15  5 */ n398;
assign n929  = /* LUT    4 11  2 */ (n21 ? n150 : n206);
assign n930  = /* LUT    9  4  7 */ (n176 ? 1'b0 : !n495);
assign n931  = /* LUT    9  7  3 */ n507;
assign n932  = /* LUT    2 14  5 */ n40;
assign n933  = /* LUT    6  7  4 */ (n131 ? (n128 ? 1'b0 : (n54 ? 1'b1 : n130)) : (n128 ? n130 : (n54 ? n130 : 1'b1)));
assign n934  = /* LUT    8  7  6 */ n438;
assign n935  = /* LUT   11  5  0 */ (n350 ? (n41 ? 1'b1 : (n6 ? 1'b1 : n92)) : 1'b0);
assign n936  = /* LUT    5  8  0 */ (n201 ? (n266 ? n193 : 1'b1) : (n266 ? (n193 ? !n270 : n270) : n270));
assign n937  = /* LUT    7  8  2 */ (n355 ? (n62 ? !n357 : 1'b1) : (n62 ? n357 : 1'b0));
assign n938  = /* LUT    7 11  7 */ (n60 ? (n59 ? n379 : n30) : n379);
assign n939  = /* LUT    5 14  7 */ n232;
assign n940  = /* LUT    6 10  5 */ (n21 ? n283 : n285);
assign n941  = /* LUT   11  9  6 */ (n105 ? !n142 : n142);
assign n942  = /* LUT    6  2  1 */ (n320 ? 1'b0 : (n322 ? 1'b0 : (n325 ? n238 : 1'b1)));
assign n943  = /* LUT    6 13  1 */ n306;
assign n944  = /* LUT    8  2  3 */ (n407 ? (n254 ? !n484 : 1'b0) : (n254 ? (n484 ? !n408 : n408) : n408));
assign n945  = /* LUT    9 11  5 */ n532;
assign n946  = /* LUT    5  6  2 */ (n205 ? (n7 ? 1'b0 : !n189) : (n7 ? (n189 ? !n201 : n201) : n201));
assign n947  = /* LUT    4 10  5 */ (n146 ? (n149 ? !n62 : 1'b1) : (n149 ? n62 : 1'b0));
assign n948  = /* LUT    6  3  2 */ (n239 ? (n87 ? n325 : (n324 ? n325 : 1'b1)) : (n87 ? 1'b0 : (n324 ? 1'b1 : n325)));
assign n949  = /* LUT    6 14  2 */ n234;
assign n950  = /* LUT    4  2  1 */ (n41 ? (n113 ? (n8 ? n42 : 1'b1) : 1'b0) : (n8 ? n42 : 1'b1));
assign n951  = /* LUT    8  3  4 */ (n415 ? (n334 ? (n46 ? n342 : 1'b1) : (n46 ? !n342 : 1'b0)) : (n334 ? (n46 ? !n342 : 1'b0) : (n46 ? n342 : 1'b1)));
assign n952  = /* LUT    7 15  0 */ n401;
assign n953  = /* LUT    5  7  3 */ (n54 ? (n130 ? n128 : (n128 ? 1'b0 : n131)) : (n130 ? n128 : (n128 ? 1'b1 : !n131)));
assign n954  = /* LUT    7  7  5 */ n143;
assign n955  = /* LUT    4  3  2 */ (n170 ? (n120 ? 1'b0 : !n117) : (n120 ? !n117 : 1'b0));
assign n956  = /* LUT    9  7  7 */ n505;
assign n957  = /* LUT    8  7  1 */ n442;
assign n958  = /* LUT    8  6  5 */ n433;
assign n959  = /* LUT    7 11  2 */ n378;
assign n960  = /* LUT    2  6  1 */ (n55 ? 1'b0 : (n49 ? 1'b0 : (n17 ? 1'b0 : !n48)));
assign n961  = /* LUT    6 10  0 */ (n21 ? !n286 : !n287);
assign n962  = /* LUT   11  9  1 */ (select ? n142 : n545);
assign n963  = /* LUT    8 10  2 */ n462;
assign n964  = /* LUT    6  2  5 */ (n327 ? (n240 ? !n326 : n326) : (n240 ? n326 : !n326));
assign n965  = /* LUT    8  2  7 */ (n412 ? n327 : !n327);
assign n966  = /* LUT    7  3  3 */ (n402 ? (n408 ? 1'b0 : !n247) : (n408 ? (n246 ? !n247 : n247) : !n246));
assign n967  = /* LUT    4 10  0 */ (n104 ? !n197 : n197);
assign n968  = /* LUT    2 10  7 */ n61;
assign n969  = /* LUT    5  6  6 */ (n180 ? (n63 ? !n127 : 1'b0) : (n63 ? (n127 ? !n144 : n144) : !n144));
assign n970  = /* LUT    6  3  6 */ (n87 ? (n239 ? (n324 ? n325 : !n325) : (n324 ? 1'b0 : n325)) : (n239 ? (n324 ? !n325 : 1'b0) : 1'b1));
assign n971  = /* LUT    6 14  6 */ n314;
assign n972  = /* LUT    4  2  5 */ (n122 ? (n123 ? 1'b0 : (n120 ? 1'b0 : !n121)) : 1'b0);
assign n973  = /* LUT   11 12  2 */ n552;
assign n974  = /* LUT   11  4  7 */ n262;
assign n975  = /* LUT    4 11  1 */ (n21 ? !n157 : !n156);
assign n976  = /* LUT    7  7  0 */ (n440 ? !n341 : n341);
assign n977  = /* LUT    9  4  6 */ (n493 ? (n424 ? (n486 ? !n420 : n420) : (n486 ? n420 : !n420)) : (n424 ? (n486 ? n420 : !n420) : (n486 ? !n420 : n420)));
assign n978  = /* LUT    5  7  7 */ (n130 ? (n131 ? (n54 ? 1'b0 : !n128) : n54) : (n131 ? (n54 ? 1'b0 : n128) : 1'b1));
assign n979  = /* LUT    9  7  2 */ n510;
assign n980  = /* LUT    4  3  6 */ (n122 ? (n123 ? 1'b0 : !n117) : (n123 ? !n117 : 1'b0));
assign n981  = /* LUT    4 14  6 */ n38;
assign n982  = /* LUT    8  6  0 */ n15;
assign n983  = /* LUT    6  9  3 */ (n21 ? n277 : n279);
assign n984  = /* LUT    5  2  4 */ (n92 ? (n116 ? 1'b0 : (n58 ? !n118 : 1'b1)) : (n58 ? !n118 : 1'b1));
assign n985  = /* LUT    4  6  7 */ !n17;
assign n986  = /* LUT    6 10  4 */ (n196 ? (n62 ? n283 : 1'b0) : (n62 ? !n283 : 1'b1));
assign n987  = /* LUT    6 13  0 */ (n304 ? (n137 ? (n282 ? !n202 : 1'b1) : (n282 ? 1'b1 : !n202)) : 1'b0);
assign n988  = /* LUT    8 10  6 */ n523;
assign n989  = /* LUT    2 10  2 */ n29;
assign n990  = /* LUT    5  6  1 */ (n189 ? (n201 ? n205 : 1'b0) : (n201 ? n7 : (n7 ? n205 : !n205)));
assign n991  = /* LUT    7  3  7 */ (n89 ? (n407 ? n247 : 1'b1) : (n246 ? (n407 ? 1'b1 : n247) : (n407 ? 1'b0 : !n247)));
assign n992  = /* LUT    4 10  4 */ (n197 ? (n62 ? !n157 : 1'b1) : (n62 ? n157 : 1'b0));
assign n993  = /* LUT    4  2  0 */ (n122 ? (n123 ? (n120 ? !n121 : 1'b0) : 1'b0) : 1'b0);
assign n994  = /* LUT    8 13  7 */ n391;
assign n995  = /* LUT   11  4  2 */ (n536 ? (n41 ? 1'b1 : (n6 ? 1'b1 : n92)) : 1'b0);
assign n996  = /* LUT    5  7  2 */ (n263 ? (n203 ? n107 : !n107) : (n203 ? !n107 : n107));
assign n999  = /* LUT    9  7  6 */ n496;
assign n1000 = /* LUT    5 13  0 */ (n227 ? (n59 ? (n60 ? !n225 : 1'b1) : 1'b1) : 1'b0);
assign n1001 = /* LUT    7 10  6 */ (n368 ? (n140 ? (n215 ? n62 : 1'b0) : (n215 ? !n62 : 1'b1)) : (n140 ? (n215 ? !n62 : 1'b1) : (n215 ? n62 : 1'b0)));
assign n1002 = /* LUT    7  2  2 */ (n87 ? (n335 ? (n323 ? !n321 : 1'b0) : (n323 ? 1'b0 : n321)) : 1'b0);
assign n1003 = /* LUT    8  6  4 */ n436;
assign n1004 = /* LUT    8  9  0 */ (n453 ? (n59 ? (n60 ? !n461 : 1'b1) : 1'b1) : 1'b0);
assign n1005 = /* LUT    6  9  7 */ (n25 ? (n62 ? n277 : 1'b0) : (n62 ? !n277 : 1'b1));
assign n1006 = /* LUT    2  6  0 */ (rst ? 1'b1 : (n44 ? n53 : 1'b0));
assign n1007 = /* LUT    5 14  1 */ n235;
assign n1008 = /* LUT    4  6  2 */ (n181 ? (n16 ? n129 : !n129) : (n16 ? !n129 : n129));
assign n1009 = /* LUT    7 14  3 */ (n60 ? (n59 ? n395 : n397) : n395);
assign n1010 = /* LUT    8 10  1 */ n465;
assign n1011 = /* LUT    6 13  4 */ n308;
assign n1012 = /* LUT    8  2  6 */ (n405 ? (n327 ? (n402 ? 1'b0 : !n89) : (n402 ? 1'b1 : n89)) : (n327 ? (n402 ? 1'b1 : n89) : (n402 ? 1'b0 : !n89)));
assign n1013 = /* LUT    7  3  2 */ (n236 ? (n331 ? (n410 ? 1'b0 : !n243) : (n410 ? 1'b1 : n243)) : (n331 ? (n410 ? 1'b1 : n243) : (n410 ? 1'b0 : !n243)));
assign n1014 = /* LUT    5  6  5 */ (n263 ? (n180 ? 1'b0 : (n178 ? n144 : !n144)) : (n180 ? (n178 ? n144 : !n144) : 1'b0));
assign n1015 = /* LUT    4  2  4 */ (n114 ? (n166 ? 1'b0 : (n118 ? 1'b1 : !n58)) : 1'b0);
assign n1016 = /* LUT    5  9  7 */ n278;
assign n1017 = /* LUT    2  5  4 */ (n95 ? !n50 : n50);
assign n1018 = /* LUT    6  5  5 */ (n50 ? (n14 ? (n51 ? 1'b1 : n52) : 1'b1) : (n14 ? 1'b1 : (n51 ? n52 : 1'b1)));
assign n1019 = /* LUT   11  4  6 */ (n56 ? (n41 ? 1'b0 : (n6 ? 1'b0 : !n92)) : 1'b0);
assign n1020 = /* LUT    8  5  7 */ n346;
assign n1021 = /* LUT    7 10  1 */ (n25 ? !n196 : n196);
assign n1022 = /* LUT    9 10  3 */ n526;
assign n1023 = /* LUT    6  9  2 */ (n204 ? n105 : !n105);
assign n1024 = /* LUT    7  2  6 */ (n335 ? n321 : !n321);
assign n1025 = /* LUT    4  9  3 */ (n197 ? (n62 ? !n148 : 1'b1) : (n62 ? n148 : 1'b0));
assign n1026 = /* LUT    8  9  4 */ n428;
assign n1027 = /* LUT    5  2  3 */ (rst ? 1'b1 : (n172 ? 1'b1 : n118));
assign n1028 = /* LUT    5 14  5 */ n86;
assign n1029 = /* LUT    4  6  6 */ (n127 ? (n184 ? (n63 ? n186 : !n186) : 1'b0) : (n184 ? 1'b0 : (n63 ? n186 : !n186)));
assign n1030 = /* LUT    7 14  7 */ n385;
assign n1031 = /* LUT    8  2  1 */ (n407 ? !n408 : 1'b0);
assign n1032 = /* LUT    6 12  3 */ n300;
assign n1033 = /* LUT    8 12  5 */ n480;
assign n1034 = /* LUT    5  6  0 */ (n107 ? (n178 ? n201 : !n201) : (n178 ? !n201 : n201));
assign n1035 = /* LUT    9  6  1 */ n502;
assign n1036 = /* LUT    2 13  3 */ n35;
assign n1037 = /* LUT    5  9  2 */ (n59 ? 1'b0 : !n60);
assign n1038 = /* LUT    4 13  5 */ (n59 ? (n60 ? n82 : n34) : n82);
assign n1039 = /* LUT    7  9  4 */ n365;
assign n1040 = /* LUT    8  5  2 */ (n430 ? (n253 ? (n414 ? !n168 : 1'b1) : (n414 ? 1'b1 : !n168)) : (n253 ? (n414 ? n168 : 1'b0) : (n414 ? 1'b0 : n168)));
assign n1041 = /* LUT    9  9  6 */ n366;
assign n1042 = /* LUT   11  3  5 */ (n254 ? !n342 : n342);
assign n1043 = /* LUT    7 10  5 */ (n368 ? (n62 ? !n369 : 1'b1) : (n62 ? n369 : 1'b0));
assign n1044 = /* LUT    7  2  1 */ (n408 ? (n402 ? 1'b0 : (n407 ? n89 : !n89)) : (n402 ? (n407 ? n89 : !n89) : 1'b0));
assign n1045 = /* LUT    8  6  3 */ (n445 ? (n346 ? n169 : 1'b1) : (n346 ? !n169 : 1'b0));
assign n1046 = /* LUT    9 10  7 */ n309;
assign n1047 = /* LUT    6  9  6 */ (n21 ? n275 : n106);
assign n1048 = /* LUT    4  6  1 */ (n127 ? !n63 : 1'b0);
assign n1049 = /* LUT    5  2  7 */ (rst ? 1'b0 : !n167);
assign n1050 = /* LUT   11  8  3 */ n454;
assign n1051 = /* LUT    8 12  0 */ n476;
assign n1052 = /* LUT    6 12  7 */ (n202 ? n307 : (n309 ? n291 : !n291));
assign n1053 = /* LUT    6  4  3 */ (n41 ? 1'b0 : !n92);
assign n1054 = /* LUT    8  4  5 */ (n409 ? 1'b0 : !n487);
assign n1055 = /* LUT    4 13  0 */ (n59 ? (n60 ? 1'b1 : !n82) : (n60 ? !n37 : 1'b1));
assign n1056 = /* LUT    8 13  1 */ (n60 ? (n59 ? n110 : n312) : n110);
assign n1057 = /* LUT    2 13  7 */ n79;
assign n1058 = /* LUT    9  6  5 */ (n503 ? (n179 ? n169 : 1'b1) : (n179 ? !n169 : 1'b0));
assign n1059 = /* LUT    5  9  6 */ (n216 ? (n263 ? !n212 : n212) : (n263 ? n212 : !n212));
assign n1060 = /* LUT    2  5  3 */ (n94 ? !n49 : n49);
assign n1061 = /* LUT    6  5  4 */ (n4 ? (n50 ? (n51 ? n260 : 1'b0) : 1'b0) : 1'b0);
assign n1062 = /* LUT    9  9  1 */ n516;
assign n1063 = /* LUT    4  5  5 */ (n25 ? n179 : !n179);
assign n1064 = /* LUT    8  5  6 */ (n349 ? (n41 ? 1'b1 : (n6 ? 1'b1 : n92)) : 1'b0);
assign n1065 = /* LUT   11 11  4 */ (n140 ? !n262 : n262);
assign n1066 = /* LUT    7 10  0 */ (n21 ? !n369 : !n371);
assign n1067 = /* LUT    5 10  7 */ n290;
assign n1068 = /* LUT    9 10  2 */ n521;
assign n1069 = /* LUT    5 13  3 */ n229;
assign n1070 = /* LUT    4  9  2 */ (n105 ? (n62 ? !n145 : 1'b1) : (n62 ? n145 : 1'b0));
assign n1071 = /* LUT    8  9  3 */ (n60 ? (n59 ? n26 : n461) : n26);
assign n1072 = /* LUT    6  8  5 */ n273;
assign n1073 = /* LUT    8  8  7 */ (n355 ? !n446 : n446);
assign n1074 = /* LUT    5  2  2 */ (n92 ? !n116 : 1'b0);
assign n1075 = /* LUT    7 13  1 */ (n390 ? (n347 ? (n367 ? !n202 : 1'b1) : (n367 ? 1'b1 : !n202)) : 1'b0);
assign n1076 = /* LUT   12  6  6 */ n553;
assign n1077 = /* LUT    5  5  4 */ n174;
assign n1078 = /* LUT    7  5  6 */ n56;
assign n1079 = /* LUT    6 12  2 */ (n60 ? (n59 ? n301 : n307) : n301);
assign n1080 = /* LUT    4 12  3 */ n90;
assign n1081 = /* LUT    8 12  4 */ n137;
assign n1082 = /* LUT    1  8  6 */ !rst;
assign n1083 = /* LUT    8  4  0 */ (n328 ? !n414 : n414);
assign n1084 = /* LUT    6  4  7 */ (n251 ? (n337 ? n245 : !n245) : (n337 ? !n245 : n245));
assign n1085 = /* LUT    9  6  0 */ n501;
assign n1086 = /* LUT    2 13  2 */ n83;
assign n1087 = /* LUT    7  6  7 */ n347;
assign n1088 = /* LUT    4 13  4 */ n161;
assign n1089 = /* LUT    7  9  3 */ (n263 ? (n7 ? (n362 ? n361 : 1'b1) : (n362 ? !n361 : 1'b0)) : (n7 ? (n362 ? !n361 : 1'b0) : (n362 ? n361 : 1'b1)));
assign n1090 = /* LUT    8 13  5 */ n481;
assign n1091 = /* LUT    8  5  1 */ (n15 ? (n41 ? 1'b0 : (n6 ? 1'b0 : !n92)) : 1'b0);
assign n1092 = /* LUT    2  5  7 */ (n98 ? !n14 : n14);
assign n1093 = /* LUT    9  9  5 */ (n513 ? (n421 ? n169 : 1'b1) : (n421 ? !n169 : 1'b0));
assign n1094 = /* LUT    6 11  6 */ (n271 ? (n62 ? !n296 : 1'b1) : (n62 ? n296 : 1'b0));
assign n1095 = /* LUT    7  2  0 */ (n410 ? !n254 : n254);
assign n1096 = /* LUT    6  8  0 */ (n25 ? (n269 ? !n197 : n197) : (n269 ? n197 : !n197));
assign n1097 = /* LUT   11  7  1 */ n542;
assign n1098 = /* LUT    8  8  2 */ n447;
assign n1099 = /* LUT   11 10  3 */ n460;
assign n1100 = /* LUT    7 13  5 */ (n389 ? (n59 ? (n60 ? !n312 : 1'b1) : 1'b1) : 1'b0);
assign n1101 = /* LUT   12  9  6 */ n543;
assign n1102 = /* LUT    9  5  3 */ (n426 ? (n12 ? 1'b0 : !n491) : (n12 ? !n492 : (n491 ? !n492 : n492)));
assign n1103 = /* LUT    6 12  6 */ n299;
assign n1104 = /* LUT    2  4  1 */ (n4 ? !n51 : 1'b0);
assign n1105 = /* LUT    6  4  2 */ (n4 ? (n91 ? !n50 : n14) : 1'b0);
assign n1106 = /* LUT    4 12  7 */ n219;
assign n1107 = /* LUT    8  4  4 */ (n488 ? (n486 ? !n420 : n420) : (n486 ? n420 : !n420));
assign n1108 = /* LUT    7  6  2 */ n309;
assign n1109 = /* LUT    9  6  4 */ n509;
assign n1110 = /* LUT    5  9  5 */ (n188 ? (n133 ? (n278 ? !n62 : 1'b1) : (n278 ? n62 : 1'b0)) : (n133 ? (n278 ? n62 : 1'b0) : (n278 ? !n62 : 1'b1)));
assign n1111 = /* LUT    9  9  0 */ n514;
assign n1112 = /* LUT    2  5  2 */ (n93 ? !n48 : n48);
assign n1113 = /* LUT    7  9  7 */ (n202 ? n461 : (n428 ? n274 : !n274));
assign n1114 = /* LUT    4  5  4 */ (select ? n179 : n125);
assign n1115 = /* LUT   11 11  3 */ (select ? n421 : n551);
assign n1116 = /* LUT    6 11  1 */ (n297 ? (n309 ? (n291 ? !n202 : 1'b1) : (n291 ? 1'b1 : !n202)) : 1'b0);
assign n1117 = /* LUT    8 11  3 */ n477;
assign n559  = /* CARRY  4  3  0 */ (n122 & 1'b0) | ((n122 | 1'b0) & n668);
assign n98   = /* CARRY  2  5  6 */ (1'b0 & n52) | ((1'b0 | n52) & n97);
assign n93   = /* CARRY  2  5  1 */ (1'b0 & n55) | ((1'b0 | n55) & n560);
assign n97   = /* CARRY  2  5  5 */ (1'b0 & n51) | ((1'b0 | n51) & n96);
assign n560  = /* CARRY  2  5  0 */ (n17 & 1'b0) | ((n17 | 1'b0) & n828);
assign n171  = /* CARRY  4  3  2 */ (1'b0 & n120) | ((1'b0 | n120) & n170);
assign n170  = /* CARRY  4  3  1 */ (1'b0 & n123) | ((1'b0 | n123) & n559);
assign n96   = /* CARRY  2  5  4 */ (1'b0 & n50) | ((1'b0 | n50) & n95);
assign n95   = /* CARRY  2  5  3 */ (1'b0 & n49) | ((1'b0 | n49) & n94);
assign n94   = /* CARRY  2  5  2 */ (1'b0 & n48) | ((1'b0 | n48) & n93);
/* FF  5 12  6 */ always @(posedge clk) if (1'b1) n221 <= 1'b0 ? 1'b0 : n561;
/* FF  9 12  1 */ always @(posedge clk) if (1'b1) n528 <= 1'b0 ? 1'b0 : n562;
/* FF  6  8  4 */ always @(posedge clk) if (1'b1) n265 <= 1'b0 ? 1'b0 : n563;
/* FF  5  4  2 */ assign n91 = n564;
/* FF  4  8  5 */ assign n104 = n565;
/* FF  7  4  4 */ assign n339 = n566;
/* FF  8  8  6 */ always @(posedge clk) if (1'b1) n450 <= 1'b0 ? 1'b0 : n567;
/* FF  7 13  0 */ assign n388 = n568;
/* FF 12  6  5 */ always @(posedge clk) if (1'b1) n554 <= 1'b0 ? 1'b0 : n569;
/* FF  5  5  3 */ always @(posedge clk) if (1'b1) n174 <= 1'b0 ? 1'b0 : n570;
/* FF  6 12  1 */ assign n84 = n571;
/* FF  7  5  5 */ assign n346 = n572;
/* FF  9  5  7 */ always @(posedge clk) if (n4) n494 <= 1'b0 ? 1'b0 : n573;
/* FF  6  4  6 */ assign n177 = n574;
/* FF  5  9  0 */ assign n201 = n575;
/* FF  7  9  2 */ assign n362 = n576;
/* FF  9  9  4 */ always @(posedge clk) if (1'b1) n70 <= 1'b0 ? 1'b0 : n577;
/* FF  5  8  4 */ assign n196 = n578;
/* FF  7  8  6 */ always @(posedge clk) if (1'b1) n359 <= 1'b0 ? 1'b0 : n579;
/* FF  2  7  6 */ always @(posedge clk) if (1'b1) n21 <= n58 ? 1'b0 : n580;
/* FF  6 11  5 */ always @(posedge clk) if (1'b1) n294 <= 1'b0 ? 1'b0 : n581;
/* FF  8 11  7 */ always @(posedge clk) if (1'b1) n473 <= 1'b0 ? 1'b0 : n582;
/* FF  5 12  1 */ assign n210 = n583;
/* FF  7 12  3 */ always @(posedge clk) if (1'b1) n382 <= 1'b0 ? 1'b0 : n584;
/* FF  4  8  0 */ assign n138 = n585;
/* FF  9 12  5 */ always @(posedge clk) if (1'b1) n530 <= 1'b0 ? 1'b0 : n586;
/* FF  2  8  7 */ always @(posedge clk) if (1'b1) n62 <= 1'b0 ? 1'b0 : n587;
/* FF  8  8  1 */ always @(posedge clk) if (1'b1) n447 <= 1'b0 ? 1'b0 : n588;
/* FF  2 11  3 */ always @(posedge clk) if (1'b1) n75 <= 1'b0 ? 1'b0 : n589;
/* FF 11 10  2 */ always @(posedge clk) if (1'b1) n547 <= 1'b0 ? 1'b0 : n590;
/* FF  7 13  4 */ assign n389 = n591;
/* FF  7  5  0 */ assign n343 = n592;
/* FF 12  9  5 */ always @(posedge clk) if (1'b1) n557 <= 1'b0 ? 1'b0 : n593;
/* FF  5  5  7 */ always @(posedge clk) if (1'b1) n175 <= 1'b0 ? 1'b0 : n594;
/* FF  9  5  2 */ assign n416 = n595;
/* FF  4 12  6 */ always @(posedge clk) if (1'b1) n160 <= 1'b0 ? 1'b0 : n596;
/* FF  8  4  3 */ assign n404 = n597;
/* FF  6 15  7 */ always @(posedge clk) if (1'b1) n319 <= 1'b0 ? 1'b0 : n598;
/* FF  6  7  3 */ assign n267 = n599;
/* FF  8  7  5 */ always @(posedge clk) if (1'b1) n441 <= 1'b0 ? 1'b0 : n600;
/* FF  7  8  1 */ assign n355 = n601;
/* FF  9  8  3 */ always @(posedge clk) if (1'b1) n509 <= n2 ? 1'b1 : n602;
/* FF  5 11  4 */ always @(posedge clk) if (1'b1) n213 <= 1'b0 ? 1'b0 : n603;
/* FF  7 11  6 */ always @(posedge clk) if (1'b1) n380 <= 1'b0 ? 1'b0 : n604;
/* FF  6 11  0 */ assign n291 = n605;
/* FF 11  9  5 */ always @(posedge clk) if (1'b1) n474 <= 1'b0 ? 1'b0 : n606;
/* FF  5 12  5 */ always @(posedge clk) if (1'b1) n220 <= 1'b0 ? 1'b0 : n607;
/* FF  9 12  0 */ always @(posedge clk) if (1'b1) n527 <= 1'b0 ? 1'b0 : n608;
/* FF  2  8  2 */ always @(posedge clk) if (1'b1) n61 <= 1'b0 ? 1'b0 : n609;
/* FF  5  4  1 */ assign n126 = n610;
/* FF  6  8  3 */ always @(posedge clk) if (1'b1) n23 <= 1'b0 ? 1'b0 : n611;
/* FF  4  8  4 */ assign n25 = n612;
/* FF  7  4  3 */ assign n10 = n613;
/* FF  8  8  5 */ always @(posedge clk) if (1'b1) n449 <= 1'b0 ? 1'b0 : n614;
/* FF  7 12  7 */ always @(posedge clk) if (1'b1) n386 <= 1'b0 ? 1'b0 : n615;
/* FF 11 10  6 */ always @(posedge clk) if (1'b1) n523 <= 1'b0 ? 1'b0 : n616;
/* FF  6  3  1 */ assign n46 = n617;
/* FF  6 14  1 */ assign n304 = n618;
/* FF  8  3  3 */ assign n413 = n619;
/* FF  6  6  6 */ always @(posedge clk) if (1'b1) n264 <= 1'b0 ? 1'b0 : n620;
/* FF  4 11  5 */ always @(posedge clk) if (1'b1) n157 <= 1'b0 ? 1'b0 : n621;
/* FF  8  7  0 */ always @(posedge clk) if (1'b1) n438 <= 1'b0 ? 1'b0 : n622;
/* FF  6  7  7 */ always @(posedge clk) if (1'b1) n143 <= n2 ? 1'b0 : n623;
/* FF 11  5  3 */ assign n12 = n624;
/* FF  5  8  3 */ assign n195 = n625;
/* FF  7 11  1 */ always @(posedge clk) if (1'b1) n377 <= 1'b0 ? 1'b0 : n626;
/* FF  4  7  7 */ assign n136 = n627;
/* FF  6 11  4 */ always @(posedge clk) if (1'b1) n290 <= 1'b0 ? 1'b0 : n628;
/* FF  8 11  6 */ always @(posedge clk) if (1'b1) n461 <= 1'b0 ? 1'b0 : n629;
/* FF  5 12  0 */ assign n216 = n630;
/* FF  5  4  5 */ assign n172 = n631;
/* FF  2 11  2 */ always @(posedge clk) if (1'b1) n30 <= 1'b0 ? 1'b0 : n632;
/* FF  7  4  7 */ assign n176 = n633;
/* FF 11 10  1 */ assign \d_out[0]  = n634;
/* FF  6  3  5 */ assign n9 = n635;
/* FF  6 14  5 */ always @(posedge clk) if (1'b1) n40 <= 1'b0 ? 1'b0 : n636;
/* FF  8  3  7 */ assign n410 = n637;
/* FF  7 15  3 */ always @(posedge clk) if (1'b1) n399 <= 1'b0 ? 1'b0 : n638;
/* FF  9  4  5 */ assign n487 = n639;
/* FF  5  7  6 */ assign n190 = n640;
/* FF  6  7  2 */ assign n144 = n641;
/* FF  8  7  4 */ always @(posedge clk) if (1'b1) n430 <= 1'b0 ? 1'b0 : n642;
/* FF 11  5  7 */ always @(posedge clk) if (1'b1) n535 <= 1'b0 ? 1'b0 : n643;
/* FF  7  8  0 */ assign n354 = n644;
/* FF  5  8  7 */ always @(posedge clk) if (1'b1) n199 <= n5 ? 1'b1 : n645;
/* FF  2  7  0 */ assign n57 = n646;
/* FF  7 11  5 */ always @(posedge clk) if (1'b1) n78 <= 1'b0 ? 1'b0 : n647;
/* FF  4  7  2 */ assign n133 = n648;
/* FF  8 11  1 */ always @(posedge clk) if (1'b1) n470 <= 1'b0 ? 1'b0 : n649;
/* FF  6 10  3 */ always @(posedge clk) if (1'b1) n285 <= 1'b0 ? 1'b0 : n650;
/* FF 11  9  4 */ always @(posedge clk) if (1'b1) n544 <= 1'b0 ? 1'b0 : n651;
/* FF  8 10  5 */ always @(posedge clk) if (1'b1) n467 <= 1'b0 ? 1'b0 : n652;
/* FF  7  4  2 */ assign n336 = n653;
/* FF  7  3  6 */ assign n333 = n654;
/* FF  4 10  3 */ always @(posedge clk) if (1'b1) n148 <= 1'b0 ? 1'b0 : n655;
/* FF  6 14  0 */ assign n311 = n656;
/* FF  6  3  0 */ assign n88 = n657;
/* FF  8  3  2 */ assign n412 = n658;
/* FF  2  2  6 */ always @(posedge clk) if (1'b1) n6 <= 1'b0 ? 1'b0 : n659;
/* FF  9  4  0 */ assign n486 = n660;
/* FF  5  7  1 */ assign n185 = n661;
/* FF  7 15  7 */ always @(posedge clk) if (1'b1) n401 <= 1'b0 ? 1'b0 : n662;
/* FF  4 11  4 */ always @(posedge clk) if (1'b1) n156 <= 1'b0 ? 1'b0 : n663;
/* FF  7  7  3 */ always @(posedge clk) if (1'b1) n90 <= 1'b0 ? 1'b0 : n664;
/* FF  6 15  1 */ always @(posedge clk) if (1'b1) n317 <= 1'b0 ? 1'b0 : n665;
/* FF  4  3  0 */ assign n666 = n667;
/* FF  9  7  5 */ always @(posedge clk) if (1'b1) n506 <= 1'b0 ? 1'b0 : n669;
/* FF  5  8  2 */ assign n194 = n670;
/* FF  7  8  4 */ always @(posedge clk) if (1'b1) n358 <= 1'b0 ? 1'b0 : n671;
/* FF  7 11  0 */ assign n376 = n672;
/* FF  9  8  6 */ always @(posedge clk) if (1'b1) n459 <= n2 ? 1'b1 : n673;
/* FF  5 11  7 */ always @(posedge clk) if (1'b1) n214 <= 1'b0 ? 1'b0 : n674;
/* FF  2  7  4 */ always @(posedge clk) if (1'b1) n59 <= n58 ? 1'b1 : n675;
/* FF  4  7  6 */ assign n135 = n676;
/* FF 11  6  3 */ always @(posedge clk) if (n4) n537 <= 1'b0 ? 1'b0 : n677;
/* FF  8 10  0 */ always @(posedge clk) if (1'b1) n462 <= 1'b0 ? 1'b0 : n678;
/* FF  6 10  7 */ always @(posedge clk) if (1'b1) n289 <= 1'b0 ? 1'b0 : n679;
/* FF  6 13  3 */ always @(posedge clk) if (1'b1) n35 <= 1'b0 ? 1'b0 : n680;
/* FF  6  2  3 */ assign n238 = n681;
/* FF  8  2  5 */ assign n248 = n682;
/* FF  7  3  1 */ assign n329 = n683;
/* FF  5  6  4 */ assign n183 = n684;
/* FF  4 10  7 */ always @(posedge clk) if (1'b1) n152 <= 1'b0 ? 1'b0 : n685;
/* FF  6  3  4 */ assign n245 = n686;
/* FF  6 14  4 */ always @(posedge clk) if (1'b1) n314 <= 1'b0 ? 1'b0 : n687;
/* FF  4  2  3 */ assign n116 = n688;
/* FF  8  3  6 */ assign n415 = n689;
/* FF  7 15  2 */ always @(posedge clk) if (1'b1) n398 <= 1'b0 ? 1'b0 : n690;
/* FF  5  7  5 */ assign n189 = n691;
/* FF  9  7  0 */ always @(posedge clk) if (1'b1) n504 <= 1'b0 ? 1'b0 : n692;
/* FF  7  7  7 */ always @(posedge clk) if (1'b1) n353 <= 1'b0 ? 1'b0 : n693;
/* FF  4  3  4 */ always @(posedge clk) if (n115) n122 <= rst ? 1'b0 : n694;
/* FF 11  5  6 */ always @(posedge clk) if (1'b1) n56 <= 1'b0 ? 1'b0 : n695;
/* FF  6  9  1 */ assign n274 = n696;
/* FF  8  6  7 */ always @(posedge clk) if (1'b1) n431 <= 1'b0 ? 1'b0 : n697;
/* FF  2  6  3 */ assign n54 = n698;
/* FF  5 14  4 */ always @(posedge clk) if (1'b1) n233 <= 1'b0 ? 1'b0 : n699;
/* FF 12  7  2 */ always @(posedge clk) if (1'b1) n556 <= 1'b0 ? 1'b0 : n700;
/* FF  6 10  2 */ always @(posedge clk) if (1'b1) n284 <= 1'b0 ? 1'b0 : n701;
/* FF  8 10  4 */ always @(posedge clk) if (1'b1) n466 <= 1'b0 ? 1'b0 : n702;
/* FF  8  2  0 */ assign n402 = n703;
/* FF  6 13  7 */ always @(posedge clk) if (1'b1) n303 <= 1'b0 ? 1'b0 : n704;
/* FF  6  2  7 */ assign n241 = n705;
/* FF  9 11  2 */ always @(posedge clk) if (1'b1) n524 <= 1'b0 ? 1'b0 : n706;
/* FF  5  3  3 */ assign n169 = n707;
/* FF  7  3  5 */ assign n332 = n708;
/* FF  4 10  2 */ always @(posedge clk) if (1'b1) n28 <= 1'b0 ? 1'b0 : n709;
/* FF  9  3  7 */ assign n342 = n710;
/* FF  8  3  1 */ assign n405 = n711;
/* FF  4  2  7 */ always @(posedge clk) if (1'b1) n41 <= 1'b0 ? 1'b0 : n712;
/* FF  5  7  0 */ assign n186 = n713;
/* FF  9  7  4 */ always @(posedge clk) if (1'b1) n489 <= 1'b0 ? 1'b0 : n714;
/* FF  5 10  2 */ always @(posedge clk) if (1'b1) n27 <= n5 ? 1'b1 : n715;
/* FF  7 10  4 */ always @(posedge clk) if (1'b1) n371 <= 1'b0 ? 1'b0 : n716;
/* FF 11  5  1 */ assign n437 = n717;
/* FF  8  6  2 */ always @(posedge clk) if (1'b1) n102 <= 1'b0 ? 1'b0 : n718;
/* FF  5 13  7 */ always @(posedge clk) if (1'b1) n231 <= 1'b0 ? 1'b0 : n719;
/* FF  2  9  4 */ always @(posedge clk) if (1'b1) n66 <= 1'b0 ? 1'b0 : n720;
/* FF  6  9  5 */ always @(posedge clk) if (1'b1) n278 <= 1'b0 ? 1'b0 : n721;
/* FF  8  9  7 */ always @(posedge clk) if (1'b1) n458 <= 1'b0 ? 1'b0 : n722;
/* FF  4  6  0 */ assign n128 = n723;
/* FF  2  6  7 */ always @(posedge clk) if (1'b1) n55 <= n1 ? 1'b0 : n724;
/* FF  5  2  6 */ always @(posedge clk) if (1'b1) n92 <= 1'b0 ? 1'b0 : n725;
/* FF  6 10  6 */ always @(posedge clk) if (1'b1) n288 <= 1'b0 ? 1'b0 : n726;
/* FF  6 13  2 */ always @(posedge clk) if (1'b1) n306 <= 1'b0 ? 1'b0 : n727;
/* FF  6  2  2 */ assign n237 = n728;
/* FF  7  3  0 */ assign n328 = n729;
/* FF  5  6  3 */ assign n63 = n730;
/* FF  4 10  6 */ always @(posedge clk) if (1'b1) n151 <= 1'b0 ? 1'b0 : n731;
/* FF  4  2  2 */ assign n115 = n732;
/* FF  8 13  0 */ always @(posedge clk) if (1'b1) n481 <= 1'b0 ? 1'b0 : n733;
/* FF  6  5  3 */ assign n257 = n734;
/* FF  8  5  5 */ assign n406 = n735;
/* FF  5 10  6 */ always @(posedge clk) if (1'b1) n207 <= n5 ? 1'b0 : n736;
/* FF  9 10  1 */ always @(posedge clk) if (1'b1) n517 <= 1'b0 ? 1'b0 : n737;
/* FF  5 13  2 */ always @(posedge clk) if (1'b1) n228 <= 1'b0 ? 1'b0 : n738;
/* FF  7  2  4 */ assign n324 = n739;
/* FF  8  6  6 */ always @(posedge clk) if (1'b1) n436 <= 1'b0 ? 1'b0 : n740;
/* FF  4  9  1 */ assign n105 = n741;
/* FF  8  9  2 */ always @(posedge clk) if (1'b1) n454 <= 1'b0 ? 1'b0 : n742;
/* FF  5 14  3 */ always @(posedge clk) if (1'b1) n232 <= 1'b0 ? 1'b0 : n743;
/* FF  6 10  1 */ always @(posedge clk) if (1'b1) n283 <= 1'b0 ? 1'b0 : n744;
/* FF  7 14  5 */ always @(posedge clk) if (1'b1) n394 <= 1'b0 ? 1'b0 : n745;
/* FF  8 10  3 */ always @(posedge clk) if (1'b1) n465 <= 1'b0 ? 1'b0 : n746;
/* FF  6  2  6 */ assign n240 = n747;
/* FF  6 13  6 */ always @(posedge clk) if (1'b1) n308 <= 1'b0 ? 1'b0 : n748;
/* FF  9 11  1 */ always @(posedge clk) if (1'b1) n498 <= 1'b0 ? 1'b0 : n749;
/* FF  7  3  4 */ assign n331 = n750;
/* FF  4 10  1 */ assign n147 = n751;
/* FF  5  6  7 */ assign n184 = n752;
/* FF  2  2  4 */ always @(posedge clk) if (1'b1) n8 <= 1'b0 ? 1'b0 : n753;
/* FF  4  2  6 */ assign n118 = n754;
/* FF  7  6  6 */ always @(posedge clk) if (n4) n350 <= 1'b0 ? 1'b0 : n755;
/* FF  4 13  3 */ always @(posedge clk) if (1'b1) n163 <= 1'b0 ? 1'b0 : n756;
/* FF  8 13  4 */ always @(posedge clk) if (1'b1) n32 <= 1'b0 ? 1'b0 : n757;
/* FF 11 12  3 */ always @(posedge clk) if (1'b1) n552 <= 1'b0 ? 1'b0 : n758;
/* FF  8  5  0 */ assign n421 = n759;
/* FF  2  5  6 */ always @(posedge clk) if (1'b1) n52 <= n1 ? 1'b0 : n760;
/* FF  6  5  7 */ always @(posedge clk) if (1'b1) n261 <= n2 ? 1'b0 : n761;
/* FF 11 11  7 */ always @(posedge clk) if (1'b1) n551 <= 1'b0 ? 1'b0 : n762;
/* FF  5 10  1 */ always @(posedge clk) if (1'b1) n206 <= n5 ? 1'b0 : n763;
/* FF  7 10  3 */ always @(posedge clk) if (1'b1) n370 <= 1'b0 ? 1'b0 : n764;
/* FF  8  6  1 */ always @(posedge clk) if (1'b1) n432 <= 1'b0 ? 1'b0 : n765;
/* FF  9 10  5 */ always @(posedge clk) if (1'b1) n521 <= 1'b0 ? 1'b0 : n766;
/* FF  5 13  6 */ always @(posedge clk) if (1'b1) n230 <= 1'b0 ? 1'b0 : n767;
/* FF  2  9  3 */ always @(posedge clk) if (1'b1) n65 <= 1'b0 ? 1'b0 : n768;
/* FF  6  9  4 */ always @(posedge clk) if (1'b1) n277 <= 1'b0 ? 1'b0 : n769;
/* FF  4  9  5 */ always @(posedge clk) if (1'b1) n72 <= 1'b0 ? 1'b0 : n770;
/* FF  8  9  6 */ always @(posedge clk) if (1'b1) n457 <= 1'b0 ? 1'b0 : n771;
/* FF 11  7  0 */ always @(posedge clk) if (1'b1) n539 <= 1'b0 ? 1'b0 : n772;
/* FF  7 14  0 */ assign n387 = n773;
/* FF  5  2  5 */ always @(posedge clk) if (1'b1) n58 <= 1'b0 ? 1'b0 : n774;
/* FF 11  8  1 */ always @(posedge clk) if (1'b1) n542 <= 1'b0 ? 1'b0 : n775;
/* FF  6 12  5 */ always @(posedge clk) if (1'b1) n300 <= 1'b0 ? 1'b0 : n776;
/* FF  6  4  1 */ assign n250 = n777;
/* FF  2 13  5 */ always @(posedge clk) if (1'b1) n82 <= 1'b0 ? 1'b0 : n778;
/* FF  5  9  4 */ assign n203 = n779;
/* FF  4 13  7 */ always @(posedge clk) if (1'b1) n34 <= 1'b0 ? 1'b0 : n780;
/* FF  6  5  2 */ assign n256 = n781;
/* FF  7  9  6 */ always @(posedge clk) if (1'b1) n365 <= 1'b0 ? 1'b0 : n782;
/* FF  2  5  1 */ assign n783 = n784;
/* FF  8  5  4 */ assign n425 = n785;
/* FF  9 10  0 */ always @(posedge clk) if (1'b1) n309 <= 1'b0 ? 1'b0 : n786;
/* FF  7 10  7 */ always @(posedge clk) if (1'b1) n373 <= 1'b0 ? 1'b0 : n787;
/* FF  5 13  1 */ assign n227 = n788;
/* FF  7  2  3 */ assign n323 = n789;
/* FF  8  9  1 */ assign n453 = n790;
/* FF  2  9  7 */ always @(posedge clk) if (1'b1) n67 <= 1'b0 ? 1'b0 : n791;
/* FF 11  7  4 */ always @(posedge clk) if (1'b1) n541 <= 1'b0 ? 1'b0 : n792;
/* FF 12  7  0 */ always @(posedge clk) if (1'b1) n555 <= 1'b0 ? 1'b0 : n793;
/* FF  4  6  3 */ assign n131 = n794;
/* FF 12  6  4 */ always @(posedge clk) if (1'b1) n553 <= 1'b0 ? 1'b0 : n795;
/* FF  5  5  2 */ assign \d_out[6]  = n796;
/* FF  7  5  4 */ assign n345 = n797;
/* FF  6 12  0 */ assign n297 = n798;
/* FF  4 12  1 */ always @(posedge clk) if (1'b1) n158 <= 1'b0 ? 1'b0 : n799;
/* FF  9  5  6 */ assign n493 = n800;
/* FF  8 12  2 */ always @(posedge clk) if (1'b1) n477 <= 1'b0 ? 1'b0 : n801;
/* FF  2  4  4 */ always @(posedge clk) if (n4) n11 <= 1'b0 ? 1'b0 : n802;
/* FF  6  4  5 */ assign n13 = n803;
/* FF  8  4  7 */ assign n262 = n804;
/* FF  2 13  0 */ always @(posedge clk) if (1'b1) n79 <= 1'b0 ? 1'b0 : n805;
/* FF  7  9  1 */ assign n281 = n806;
/* FF  9  6  7 */ always @(posedge clk) if (1'b1) n503 <= 1'b0 ? 1'b0 : n807;
/* FF  9  9  3 */ always @(posedge clk) if (1'b1) n514 <= 1'b0 ? 1'b0 : n808;
/* FF  2  5  5 */ always @(posedge clk) if (1'b1) n51 <= n1 ? 1'b0 : n809;
/* FF  6  5  6 */ assign n260 = n810;
/* FF  7 10  2 */ always @(posedge clk) if (1'b1) n369 <= 1'b0 ? 1'b0 : n811;
/* FF  9 10  4 */ always @(posedge clk) if (1'b1) n520 <= 1'b0 ? 1'b0 : n812;
/* FF  5 13  5 */ always @(posedge clk) if (1'b1) n229 <= 1'b0 ? 1'b0 : n813;
/* FF  2  9  2 */ assign n64 = n814;
/* FF  7  2  7 */ assign n326 = n815;
/* FF  4  9  4 */ always @(posedge clk) if (1'b1) n71 <= 1'b0 ? 1'b0 : n816;
/* FF  8  8  0 */ assign n446 = n817;
/* FF  6  8  7 */ always @(posedge clk) if (1'b1) n273 <= 1'b0 ? 1'b0 : n818;
/* FF  9 13  5 */ always @(posedge clk) if (1'b1) n532 <= n2 ? 1'b1 : n819;
/* FF  9  5  1 */ assign n490 = n820;
/* FF  6  4  0 */ assign n249 = n821;
/* FF  8 12  6 */ always @(posedge clk) if (1'b1) n480 <= 1'b0 ? 1'b0 : n822;
/* FF  8  4  2 */ assign n418 = n823;
/* FF  9  6  2 */ always @(posedge clk) if (1'b1) n137 <= 1'b0 ? 1'b0 : n824;
/* FF  2 13  4 */ always @(posedge clk) if (1'b1) n38 <= 1'b0 ? 1'b0 : n825;
/* FF  2  5  0 */ assign n826 = n827;
/* FF  4 13  6 */ always @(posedge clk) if (1'b1) n165 <= 1'b0 ? 1'b0 : n829;
/* FF  6  5  1 */ assign n255 = n830;
/* FF  7  9  5 */ always @(posedge clk) if (1'b1) n364 <= 1'b0 ? 1'b0 : n831;
/* FF 11 11  1 */ assign \d_out[1]  = n832;
/* FF  8  5  3 */ assign n424 = n833;
/* FF  9  9  7 */ always @(posedge clk) if (1'b1) n497 <= 1'b0 ? 1'b0 : n834;
/* FF  5 12  4 */ always @(posedge clk) if (1'b1) n219 <= 1'b0 ? 1'b0 : n835;
/* FF  7 12  6 */ always @(posedge clk) if (1'b1) n385 <= 1'b0 ? 1'b0 : n836;
/* FF 11  7  3 */ always @(posedge clk) if (1'b1) n540 <= 1'b0 ? 1'b0 : n837;
/* FF  4  8  3 */ assign n140 = n838;
/* FF  2 11  6 */ always @(posedge clk) if (1'b1) n77 <= 1'b0 ? 1'b0 : n839;
/* FF  7 13  7 */ always @(posedge clk) if (1'b1) n391 <= 1'b0 ? 1'b0 : n840;
/* FF  7  5  3 */ assign n344 = n841;
/* FF  9  5  5 */ assign n492 = n842;
/* FF  2 12  7 */ always @(posedge clk) if (1'b1) n31 <= 1'b0 ? 1'b0 : n843;
/* FF  8 12  1 */ always @(posedge clk) if (1'b1) n476 <= 1'b0 ? 1'b0 : n844;
/* FF  2  4  3 */ assign n45 = n845;
/* FF  6  4  4 */ assign n252 = n846;
/* FF  8  4  6 */ assign n420 = n847;
/* FF  6  7  6 */ assign n270 = n848;
/* FF  7  9  0 */ assign n361 = n849;
/* FF  9  9  2 */ always @(posedge clk) if (1'b1) n513 <= 1'b0 ? 1'b0 : n850;
/* FF  6 11  3 */ always @(posedge clk) if (1'b1) n293 <= 1'b0 ? 1'b0 : n851;
/* FF  7 12  1 */ always @(posedge clk) if (1'b1) n109 <= 1'b0 ? 1'b0 : n852;
/* FF  9 12  3 */ always @(posedge clk) if (1'b1) n529 <= 1'b0 ? 1'b0 : n853;
/* FF  6  8  6 */ always @(posedge clk) if (1'b1) n272 <= 1'b0 ? 1'b0 : n854;
/* FF  2 11  1 */ always @(posedge clk) if (1'b1) n74 <= 1'b0 ? 1'b0 : n855;
/* FF  7  4  6 */ assign n341 = n856;
/* FF  4  8  7 */ assign n141 = n857;
/* FF  7  5  7 */ always @(posedge clk) if (1'b1) n348 <= 1'b0 ? 1'b0 : n858;
/* FF  4 12  4 */ always @(posedge clk) if (1'b1) n85 <= 1'b0 ? 1'b0 : n859;
/* FF  8  4  1 */ assign n408 = n860;
/* FF  6 15  5 */ always @(posedge clk) if (1'b1) n310 <= 1'b0 ? 1'b0 : n861;
/* FF  6  7  1 */ assign n266 = n862;
/* FF  8  7  3 */ always @(posedge clk) if (1'b1) n440 <= 1'b0 ? 1'b0 : n863;
/* FF  5  8  6 */ assign n198 = n864;
/* FF  9  8  1 */ assign \d_out[3]  = n865;
/* FF  5 11  2 */ assign n212 = n866;
/* FF  7 11  4 */ always @(posedge clk) if (1'b1) n379 <= 1'b0 ? 1'b0 : n867;
/* FF  4  7  1 */ assign n20 = n868;
/* FF  8 11  0 */ always @(posedge clk) if (1'b1) n469 <= 1'b0 ? 1'b0 : n869;
/* FF  6 11  7 */ always @(posedge clk) if (1'b1) n296 <= 1'b0 ? 1'b0 : n870;
/* FF 11  9  3 */ always @(posedge clk) if (1'b1) n543 <= 1'b0 ? 1'b0 : n871;
/* FF  5 12  3 */ always @(posedge clk) if (1'b1) n218 <= 1'b0 ? 1'b0 : n872;
/* FF  7 12  5 */ always @(posedge clk) if (1'b1) n384 <= 1'b0 ? 1'b0 : n873;
/* FF  4  8  2 */ assign n139 = n874;
/* FF  7  4  1 */ assign n338 = n875;
/* FF  2 11  5 */ always @(posedge clk) if (1'b1) n76 <= 1'b0 ? 1'b0 : n876;
/* FF 11 10  4 */ always @(posedge clk) if (1'b1) n526 <= 1'b0 ? 1'b0 : n877;
/* FF  7  5  2 */ assign n179 = n878;
/* FF  9  5  4 */ assign n491 = n879;
/* FF  2  4  2 */ assign n44 = n880;
/* FF  4 11  3 */ always @(posedge clk) if (1'b1) n155 <= 1'b0 ? 1'b0 : n881;
/* FF  6 15  0 */ always @(posedge clk) if (1'b1) n316 <= 1'b0 ? 1'b0 : n882;
/* FF  6  7  5 */ assign n269 = n883;
/* FF 11 13  5 */ always @(posedge clk) if (1'b1) n110 <= 1'b0 ? 1'b0 : n884;
/* FF  8  7  7 */ always @(posedge clk) if (1'b1) n443 <= 1'b0 ? 1'b0 : n885;
/* FF  5  8  1 */ assign n193 = n886;
/* FF  7  8  3 */ always @(posedge clk) if (1'b1) n357 <= 1'b0 ? 1'b0 : n887;
/* FF  9  8  5 */ always @(posedge clk) if (1'b1) n510 <= n2 ? 1'b1 : n888;
/* FF  5 11  6 */ always @(posedge clk) if (1'b1) n108 <= 1'b0 ? 1'b0 : n889;
/* FF  4  7  5 */ assign n134 = n890;
/* FF  6 11  2 */ always @(posedge clk) if (1'b1) n292 <= 1'b0 ? 1'b0 : n891;
/* FF 11  6  2 */ always @(posedge clk) if (n4) n536 <= 1'b0 ? 1'b0 : n892;
/* FF  8 11  4 */ always @(posedge clk) if (1'b1) n472 <= 1'b0 ? 1'b0 : n893;
/* FF 11  9  7 */ always @(posedge clk) if (1'b1) n26 <= 1'b0 ? 1'b0 : n894;
/* FF  7 12  0 */ assign n211 = n895;
/* FF  5 12  7 */ always @(posedge clk) if (1'b1) n222 <= 1'b0 ? 1'b0 : n896;
/* FF  4  8  6 */ assign n22 = n897;
/* FF  7  4  5 */ assign n340 = n898;
/* FF  2 11  0 */ always @(posedge clk) if (1'b1) n73 <= 1'b0 ? 1'b0 : n899;
/* FF  6 14  3 */ always @(posedge clk) if (1'b1) n313 <= 1'b0 ? 1'b0 : n900;
/* FF  6  3  3 */ assign n244 = n901;
/* FF  8  3  5 */ assign n407 = n902;
/* FF 12  9  2 */ always @(posedge clk) if (1'b1) n374 <= 1'b0 ? 1'b0 : n903;
/* FF  7 15  1 */ always @(posedge clk) if (1'b1) n397 <= 1'b0 ? 1'b0 : n904;
/* FF  9  4  3 */ assign n484 = n905;
/* FF  5  7  4 */ assign n188 = n906;
/* FF  6 15  4 */ always @(posedge clk) if (1'b1) n318 <= 1'b0 ? 1'b0 : n907;
/* FF  4  3  3 */ always @(posedge clk) if (n115) n121 <= rst ? 1'b0 : n908;
/* FF  6  7  0 */ assign n200 = n909;
/* FF  8  7  2 */ always @(posedge clk) if (1'b1) n429 <= 1'b0 ? 1'b0 : n910;
/* FF 11  5  5 */ always @(posedge clk) if (1'b1) n99 <= 1'b0 ? 1'b0 : n911;
/* FF  5  8  5 */ assign n197 = n912;
/* FF  9  8  0 */ assign n2 = n913;
/* FF  7  8  7 */ always @(posedge clk) if (1'b1) n360 <= 1'b0 ? 1'b0 : n914;
/* FF  5 11  1 */ assign n178 = n915;
/* FF  7 11  3 */ always @(posedge clk) if (1'b1) n378 <= 1'b0 ? 1'b0 : n916;
/* FF  4  7  0 */ assign n132 = n917;
/* FF  2  7  7 */ always @(posedge clk) if (1'b1) n60 <= n58 ? 1'b1 : n918;
/* FF 11  6  6 */ always @(posedge clk) if (n4) n538 <= 1'b0 ? 1'b0 : n919;
/* FF  5 12  2 */ always @(posedge clk) if (1'b1) n217 <= 1'b0 ? 1'b0 : n920;
/* FF  7 12  4 */ always @(posedge clk) if (1'b1) n383 <= 1'b0 ? 1'b0 : n921;
/* FF  4  8  1 */ assign n5 = n922;
/* FF  7  4  0 */ assign n337 = n923;
/* FF  9 12  6 */ always @(posedge clk) if (1'b1) n531 <= 1'b0 ? 1'b0 : n924;
/* FF  8  3  0 */ assign n411 = n925;
/* FF  6  3  7 */ assign n247 = n926;
/* FF  6  6  3 */ assign \d_out[5]  = n927;
/* FF  7 15  5 */ always @(posedge clk) if (1'b1) n400 <= 1'b0 ? 1'b0 : n928;
/* FF  4 11  2 */ always @(posedge clk) if (1'b1) n154 <= 1'b0 ? 1'b0 : n929;
/* FF  9  4  7 */ assign n485 = n930;
/* FF  9  7  3 */ always @(posedge clk) if (1'b1) n392 <= 1'b0 ? 1'b0 : n931;
/* FF  2 14  5 */ always @(posedge clk) if (1'b1) n86 <= 1'b0 ? 1'b0 : n932;
/* FF  6  7  4 */ assign n268 = n933;
/* FF  8  7  6 */ always @(posedge clk) if (1'b1) n442 <= 1'b0 ? 1'b0 : n934;
/* FF 11  5  0 */ assign n499 = n935;
/* FF  5  8  0 */ assign n192 = n936;
/* FF  7  8  2 */ always @(posedge clk) if (1'b1) n356 <= 1'b0 ? 1'b0 : n937;
/* FF  7 11  7 */ always @(posedge clk) if (1'b1) n381 <= 1'b0 ? 1'b0 : n938;
/* FF  5 14  7 */ always @(posedge clk) if (1'b1) n235 <= 1'b0 ? 1'b0 : n939;
/* FF  6 10  5 */ always @(posedge clk) if (1'b1) n287 <= 1'b0 ? 1'b0 : n940;
/* FF 11  9  6 */ always @(posedge clk) if (1'b1) n545 <= 1'b0 ? 1'b0 : n941;
/* FF  6  2  1 */ assign n236 = n942;
/* FF  6 13  1 */ always @(posedge clk) if (1'b1) n305 <= 1'b0 ? 1'b0 : n943;
/* FF  8  2  3 */ assign n403 = n944;
/* FF  9 11  5 */ always @(posedge clk) if (1'b1) n525 <= 1'b0 ? 1'b0 : n945;
/* FF  5  6  2 */ assign n182 = n946;
/* FF  4 10  5 */ always @(posedge clk) if (1'b1) n150 <= 1'b0 ? 1'b0 : n947;
/* FF  6  3  2 */ assign n243 = n948;
/* FF  6 14  2 */ always @(posedge clk) if (1'b1) n312 <= 1'b0 ? 1'b0 : n949;
/* FF  4  2  1 */ assign n114 = n950;
/* FF  8  3  4 */ assign n414 = n951;
/* FF  7 15  0 */ always @(posedge clk) if (1'b1) n396 <= 1'b0 ? 1'b0 : n952;
/* FF  5  7  3 */ assign n187 = n953;
/* FF  7  7  5 */ always @(posedge clk) if (1'b1) n352 <= 1'b0 ? 1'b0 : n954;
/* FF  4  3  2 */ always @(posedge clk) if (n115) n120 <= rst ? 1'b0 : n955;
/* FF  9  7  7 */ always @(posedge clk) if (1'b1) n507 <= 1'b0 ? 1'b0 : n956;
/* FF  8  7  1 */ always @(posedge clk) if (1'b1) n439 <= 1'b0 ? 1'b0 : n957;
/* FF  8  6  5 */ always @(posedge clk) if (1'b1) n435 <= 1'b0 ? 1'b0 : n958;
/* FF  7 11  2 */ always @(posedge clk) if (1'b1) n224 <= 1'b0 ? 1'b0 : n959;
/* FF  2  6  1 */ assign n53 = n960;
/* FF  6 10  0 */ assign n282 = n961;
/* FF 11  9  1 */ assign \d_out[4]  = n962;
/* FF  8 10  2 */ always @(posedge clk) if (1'b1) n464 <= 1'b0 ? 1'b0 : n963;
/* FF  6  2  5 */ assign n239 = n964;
/* FF  8  2  7 */ assign n335 = n965;
/* FF  7  3  3 */ assign n173 = n966;
/* FF  4 10  0 */ assign n146 = n967;
/* FF  2 10  7 */ always @(posedge clk) if (1'b1) n69 <= n5 ? 1'b1 : n968;
/* FF  5  6  6 */ assign n101 = n969;
/* FF  6  3  6 */ assign n246 = n970;
/* FF  6 14  6 */ always @(posedge clk) if (1'b1) n315 <= 1'b0 ? 1'b0 : n971;
/* FF  4  2  5 */ assign n42 = n972;
/* FF 11 12  2 */ always @(posedge clk) if (1'b1) n533 <= 1'b0 ? 1'b0 : n973;
/* FF 11  4  7 */ always @(posedge clk) if (1'b1) n534 <= n2 ? 1'b1 : n974;
/* FF  4 11  1 */ assign n153 = n975;
/* FF  7  7  0 */ assign n142 = n976;
/* FF  9  4  6 */ assign n254 = n977;
/* FF  5  7  7 */ assign n191 = n978;
/* FF  9  7  2 */ always @(posedge clk) if (1'b1) n505 <= 1'b0 ? 1'b0 : n979;
/* FF  4  3  6 */ always @(posedge clk) if (n115) n123 <= rst ? 1'b0 : n980;
/* FF  4 14  6 */ always @(posedge clk) if (1'b1) n111 <= 1'b0 ? 1'b0 : n981;
/* FF  8  6  0 */ always @(posedge clk) if (1'b1) n428 <= 1'b0 ? 1'b0 : n982;
/* FF  6  9  3 */ always @(posedge clk) if (1'b1) n276 <= 1'b0 ? 1'b0 : n983;
/* FF  5  2  4 */ assign n167 = n984;
/* FF  4  6  7 */ always @(posedge clk) if (1'b1) n17 <= n1 ? 1'b0 : n985;
/* FF  6 10  4 */ always @(posedge clk) if (1'b1) n286 <= 1'b0 ? 1'b0 : n986;
/* FF  6 13  0 */ assign n263 = n987;
/* FF  8 10  6 */ always @(posedge clk) if (1'b1) n468 <= 1'b0 ? 1'b0 : n988;
/* FF  2 10  2 */ always @(posedge clk) if (1'b1) n68 <= n5 ? 1'b0 : n989;
/* FF  5  6  1 */ assign n181 = n990;
/* FF  7  3  7 */ assign n334 = n991;
/* FF  4 10  4 */ always @(posedge clk) if (1'b1) n149 <= 1'b0 ? 1'b0 : n992;
/* FF  4  2  0 */ assign n113 = n993;
/* FF  8 13  7 */ always @(posedge clk) if (1'b1) n483 <= 1'b0 ? 1'b0 : n994;
/* FF 11  4  2 */ assign n409 = n995;
/* FF  5  7  2 */ assign n127 = n996;
/* FF  4  3  1 */ assign n997 = n998;
/* FF  9  7  6 */ always @(posedge clk) if (1'b1) n460 <= 1'b0 ? 1'b0 : n999;
/* FF  5 13  0 */ assign n226 = n1000;
/* FF  7 10  6 */ always @(posedge clk) if (1'b1) n372 <= 1'b0 ? 1'b0 : n1001;
/* FF  7  2  2 */ assign n322 = n1002;
/* FF  8  6  4 */ always @(posedge clk) if (1'b1) n434 <= 1'b0 ? 1'b0 : n1003;
/* FF  8  9  0 */ assign n452 = n1004;
/* FF  6  9  7 */ always @(posedge clk) if (1'b1) n280 <= 1'b0 ? 1'b0 : n1005;
/* FF  2  6  0 */ assign n47 = n1006;
/* FF  5 14  1 */ always @(posedge clk) if (1'b1) n225 <= 1'b0 ? 1'b0 : n1007;
/* FF  4  6  2 */ assign n130 = n1008;
/* FF  7 14  3 */ always @(posedge clk) if (1'b1) n393 <= 1'b0 ? 1'b0 : n1009;
/* FF  8 10  1 */ always @(posedge clk) if (1'b1) n463 <= 1'b0 ? 1'b0 : n1010;
/* FF  6 13  4 */ always @(posedge clk) if (1'b1) n307 <= 1'b0 ? 1'b0 : n1011;
/* FF  8  2  6 */ assign n87 = n1012;
/* FF  7  3  2 */ assign n330 = n1013;
/* FF  5  6  5 */ assign n18 = n1014;
/* FF  4  2  4 */ assign n117 = n1015;
/* FF  5  9  7 */ always @(posedge clk) if (1'b1) n106 <= n5 ? 1'b0 : n1016;
/* FF  2  5  4 */ always @(posedge clk) if (1'b1) n50 <= n1 ? 1'b0 : n1017;
/* FF  6  5  5 */ assign n259 = n1018;
/* FF 11  4  6 */ assign n495 = n1019;
/* FF  8  5  7 */ always @(posedge clk) if (1'b1) n427 <= n2 ? 1'b0 : n1020;
/* FF  7 10  1 */ assign n368 = n1021;
/* FF  9 10  3 */ always @(posedge clk) if (1'b1) n519 <= 1'b0 ? 1'b0 : n1022;
/* FF  6  9  2 */ always @(posedge clk) if (1'b1) n275 <= 1'b0 ? 1'b0 : n1023;
/* FF  7  2  6 */ assign n325 = n1024;
/* FF  4  9  3 */ always @(posedge clk) if (1'b1) n145 <= 1'b0 ? 1'b0 : n1025;
/* FF  8  9  4 */ always @(posedge clk) if (1'b1) n456 <= 1'b0 ? 1'b0 : n1026;
/* FF  5  2  3 */ assign n1 = n1027;
/* FF  5 14  5 */ always @(posedge clk) if (1'b1) n234 <= 1'b0 ? 1'b0 : n1028;
/* FF  4  6  6 */ assign n16 = n1029;
/* FF  7 14  7 */ always @(posedge clk) if (1'b1) n395 <= 1'b0 ? 1'b0 : n1030;
/* FF  8  2  1 */ assign n327 = n1031;
/* FF  6 12  3 */ always @(posedge clk) if (1'b1) n299 <= 1'b0 ? 1'b0 : n1032;
/* FF  8 12  5 */ always @(posedge clk) if (1'b1) n479 <= 1'b0 ? 1'b0 : n1033;
/* FF  5  6  0 */ assign n180 = n1034;
/* FF  9  6  1 */ always @(posedge clk) if (1'b1) n444 <= 1'b0 ? 1'b0 : n1035;
/* FF  2 13  3 */ always @(posedge clk) if (1'b1) n81 <= 1'b0 ? 1'b0 : n1036;
/* FF  5  9  2 */ assign n202 = n1037;
/* FF  4 13  5 */ always @(posedge clk) if (1'b1) n164 <= 1'b0 ? 1'b0 : n1038;
/* FF  7  9  4 */ always @(posedge clk) if (1'b1) n363 <= 1'b0 ? 1'b0 : n1039;
/* FF  8  5  2 */ assign n423 = n1040;
/* FF  9  9  6 */ always @(posedge clk) if (1'b1) n516 <= 1'b0 ? 1'b0 : n1041;
/* FF 11  3  5 */ assign n89 = n1042;
/* FF  7 10  5 */ always @(posedge clk) if (1'b1) n215 <= 1'b0 ? 1'b0 : n1043;
/* FF  7  2  1 */ assign n321 = n1044;
/* FF  8  6  3 */ always @(posedge clk) if (1'b1) n433 <= 1'b0 ? 1'b0 : n1045;
/* FF  9 10  7 */ always @(posedge clk) if (1'b1) n522 <= 1'b0 ? 1'b0 : n1046;
/* FF  6  9  6 */ always @(posedge clk) if (1'b1) n279 <= 1'b0 ? 1'b0 : n1047;
/* FF  4  6  1 */ assign n129 = n1048;
/* FF  5  2  7 */ always @(posedge clk) if (1'b1) n4 <= 1'b0 ? 1'b0 : n1049;
/* FF 11  8  3 */ always @(posedge clk) if (1'b1) n511 <= 1'b0 ? 1'b0 : n1050;
/* FF  8 12  0 */ always @(posedge clk) if (1'b1) n475 <= 1'b0 ? 1'b0 : n1051;
/* FF  6 12  7 */ always @(posedge clk) if (1'b1) n302 <= 1'b0 ? 1'b0 : n1052;
/* FF  6  4  3 */ assign n168 = n1053;
/* FF  8  4  5 */ assign n242 = n1054;
/* FF  4 13  0 */ assign n162 = n1055;
/* FF  8 13  1 */ always @(posedge clk) if (1'b1) n482 <= 1'b0 ? 1'b0 : n1056;
/* FF  2 13  7 */ always @(posedge clk) if (1'b1) n83 <= 1'b0 ? 1'b0 : n1057;
/* FF  9  6  5 */ always @(posedge clk) if (1'b1) n502 <= 1'b0 ? 1'b0 : n1058;
/* FF  5  9  6 */ assign n205 = n1059;
/* FF  2  5  3 */ always @(posedge clk) if (1'b1) n49 <= n1 ? 1'b0 : n1060;
/* FF  6  5  4 */ assign n258 = n1061;
/* FF  9  9  1 */ always @(posedge clk) if (1'b1) n209 <= 1'b0 ? 1'b0 : n1062;
/* FF  4  5  5 */ always @(posedge clk) if (1'b1) n125 <= 1'b0 ? 1'b0 : n1063;
/* FF  8  5  6 */ assign n426 = n1064;
/* FF 11 11  4 */ always @(posedge clk) if (1'b1) n550 <= 1'b0 ? 1'b0 : n1065;
/* FF  7 10  0 */ assign n367 = n1066;
/* FF  5 10  7 */ always @(posedge clk) if (1'b1) n208 <= n5 ? 1'b0 : n1067;
/* FF  9 10  2 */ always @(posedge clk) if (1'b1) n518 <= 1'b0 ? 1'b0 : n1068;
/* FF  5 13  3 */ always @(posedge clk) if (1'b1) n36 <= 1'b0 ? 1'b0 : n1069;
/* FF  4  9  2 */ always @(posedge clk) if (1'b1) n29 <= 1'b0 ? 1'b0 : n1070;
/* FF  8  9  3 */ always @(posedge clk) if (1'b1) n455 <= 1'b0 ? 1'b0 : n1071;
/* FF  6  8  5 */ always @(posedge clk) if (1'b1) n24 <= 1'b0 ? 1'b0 : n1072;
/* FF  8  8  7 */ always @(posedge clk) if (1'b1) n451 <= 1'b0 ? 1'b0 : n1073;
/* FF  5  2  2 */ assign n166 = n1074;
/* FF  7 13  1 */ assign n7 = n1075;
/* FF 12  6  6 */ always @(posedge clk) if (1'b1) n445 <= 1'b0 ? 1'b0 : n1076;
/* FF  5  5  4 */ always @(posedge clk) if (1'b1) n15 <= 1'b0 ? 1'b0 : n1077;
/* FF  7  5  6 */ always @(posedge clk) if (1'b1) n347 <= 1'b0 ? 1'b0 : n1078;
/* FF  6 12  2 */ always @(posedge clk) if (1'b1) n298 <= 1'b0 ? 1'b0 : n1079;
/* FF  4 12  3 */ always @(posedge clk) if (1'b1) n159 <= 1'b0 ? 1'b0 : n1080;
/* FF  8 12  4 */ always @(posedge clk) if (1'b1) n478 <= 1'b0 ? 1'b0 : n1081;
/* FF  1  8  6 */ always @(posedge clk) if (n47) d_vld <= 1'b0 ? 1'b0 : n1082;
/* FF  8  4  0 */ assign n417 = n1083;
/* FF  6  4  7 */ assign n253 = n1084;
/* FF  9  6  0 */ always @(posedge clk) if (1'b1) n500 <= 1'b0 ? 1'b0 : n1085;
/* FF  2 13  2 */ always @(posedge clk) if (1'b1) n80 <= 1'b0 ? 1'b0 : n1086;
/* FF  7  6  7 */ always @(posedge clk) if (n4) n351 <= 1'b0 ? 1'b0 : n1087;
/* FF  4 13  4 */ always @(posedge clk) if (1'b1) n37 <= 1'b0 ? 1'b0 : n1088;
/* FF  7  9  3 */ assign n107 = n1089;
/* FF  8 13  5 */ always @(posedge clk) if (1'b1) n33 <= 1'b0 ? 1'b0 : n1090;
/* FF  8  5  1 */ assign n422 = n1091;
/* FF  2  5  7 */ always @(posedge clk) if (1'b1) n14 <= n1 ? 1'b0 : n1092;
/* FF  9  9  5 */ always @(posedge clk) if (1'b1) n515 <= 1'b0 ? 1'b0 : n1093;
/* FF  6 11  6 */ always @(posedge clk) if (1'b1) n295 <= 1'b0 ? 1'b0 : n1094;
/* FF  7  2  0 */ assign n320 = n1095;
/* FF  6  8  0 */ assign n271 = n1096;
/* FF 11  7  1 */ always @(posedge clk) if (1'b1) n496 <= 1'b0 ? 1'b0 : n1097;
/* FF  8  8  2 */ always @(posedge clk) if (1'b1) n448 <= 1'b0 ? 1'b0 : n1098;
/* FF 11 10  3 */ always @(posedge clk) if (1'b1) n548 <= 1'b0 ? 1'b0 : n1099;
/* FF  7 13  5 */ assign n390 = n1100;
/* FF 12  9  6 */ always @(posedge clk) if (1'b1) n558 <= 1'b0 ? 1'b0 : n1101;
/* FF  9  5  3 */ assign n488 = n1102;
/* FF  6 12  6 */ always @(posedge clk) if (1'b1) n301 <= 1'b0 ? 1'b0 : n1103;
/* FF  2  4  1 */ assign n43 = n1104;
/* FF  6  4  2 */ assign n251 = n1105;
/* FF  4 12  7 */ always @(posedge clk) if (1'b1) n161 <= 1'b0 ? 1'b0 : n1106;
/* FF  8  4  4 */ assign n419 = n1107;
/* FF  7  6  2 */ always @(posedge clk) if (n4) n349 <= 1'b0 ? 1'b0 : n1108;
/* FF  9  6  4 */ always @(posedge clk) if (1'b1) n501 <= 1'b0 ? 1'b0 : n1109;
/* FF  5  9  5 */ assign n204 = n1110;
/* FF  9  9  0 */ always @(posedge clk) if (1'b1) n512 <= 1'b0 ? 1'b0 : n1111;
/* FF  2  5  2 */ always @(posedge clk) if (1'b1) n48 <= n1 ? 1'b0 : n1112;
/* FF  7  9  7 */ always @(posedge clk) if (1'b1) n366 <= 1'b0 ? 1'b0 : n1113;
/* FF  4  5  4 */ assign \d_out[7]  = n1114;
/* FF 11 11  3 */ assign \d_out[2]  = n1115;
/* FF  6 11  1 */ assign n103 = n1116;
/* FF  8 11  3 */ always @(posedge clk) if (1'b1) n471 <= 1'b0 ? 1'b0 : n1117;

endmodule

