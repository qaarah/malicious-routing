module top (input a, b, output y);

assign y = a & b;
//  assign y = (s)?b:(a & b);

endmodule
